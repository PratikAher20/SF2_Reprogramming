`timescale 1 ns/100 ps
// Version: v11.8 11.8.0.26


module TAMPER(
       JTAG_ACTIVE,
       LOCK_TAMPER_DETECT,
       MESH_SHORT_ERROR,
       CLK_ERROR,
       DETECT_CATEGORY,
       DETECT_ATTEMPT,
       DETECT_FAIL,
       DIGEST_ERROR,
       POWERUP_DIGEST_ERROR,
       SC_ROM_DIGEST_ERROR,
       TAMPER_CHANGE_STROBE,
       LOCKDOWN_ALL_N,
       DISABLE_ALL_IOS_N,
       RESET_N,
       ZEROIZE_N
    );
output JTAG_ACTIVE;
output LOCK_TAMPER_DETECT;
output MESH_SHORT_ERROR;
output CLK_ERROR;
output [3:0] DETECT_CATEGORY;
output DETECT_ATTEMPT;
output DETECT_FAIL;
output DIGEST_ERROR;
output POWERUP_DIGEST_ERROR;
output SC_ROM_DIGEST_ERROR;
output TAMPER_CHANGE_STROBE;
input  LOCKDOWN_ALL_N;
input  DISABLE_ALL_IOS_N;
input  RESET_N;
input  ZEROIZE_N;

    parameter ZEROIZE_CONFIG = "" ;
    parameter POWERUP_DIGEST_ERROR_CONFIG = "" ;
    parameter CLK_ERROR_CONFIG = 0 ;
    
endmodule


module RCOSC_25_50MHZ(
       CLKOUT
    );
output CLKOUT;

    parameter FREQUENCY = 50.0 ;
    
endmodule


module MSS_075(
       CAN_RXBUS_MGPIO3A_H2F_A,
       CAN_RXBUS_MGPIO3A_H2F_B,
       CAN_TX_EBL_MGPIO4A_H2F_A,
       CAN_TX_EBL_MGPIO4A_H2F_B,
       CAN_TXBUS_MGPIO2A_H2F_A,
       CAN_TXBUS_MGPIO2A_H2F_B,
       CLK_CONFIG_APB,
       COMMS_INT,
       CONFIG_PRESET_N,
       EDAC_ERROR,
       F_FM0_RDATA,
       F_FM0_READYOUT,
       F_FM0_RESP,
       F_HM0_ADDR,
       F_HM0_ENABLE,
       F_HM0_SEL,
       F_HM0_SIZE,
       F_HM0_TRANS1,
       F_HM0_WDATA,
       F_HM0_WRITE,
       FAB_CHRGVBUS,
       FAB_DISCHRGVBUS,
       FAB_DMPULLDOWN,
       FAB_DPPULLDOWN,
       FAB_DRVVBUS,
       FAB_IDPULLUP,
       FAB_OPMODE,
       FAB_SUSPENDM,
       FAB_TERMSEL,
       FAB_TXVALID,
       FAB_VCONTROL,
       FAB_VCONTROLLOADM,
       FAB_XCVRSEL,
       FAB_XDATAOUT,
       FACC_GLMUX_SEL,
       FIC32_0_MASTER,
       FIC32_1_MASTER,
       FPGA_RESET_N,
       GTX_CLK,
       H2F_INTERRUPT,
       H2F_NMI,
       H2FCALIB,
       I2C0_SCL_MGPIO31B_H2F_A,
       I2C0_SCL_MGPIO31B_H2F_B,
       I2C0_SDA_MGPIO30B_H2F_A,
       I2C0_SDA_MGPIO30B_H2F_B,
       I2C1_SCL_MGPIO1A_H2F_A,
       I2C1_SCL_MGPIO1A_H2F_B,
       I2C1_SDA_MGPIO0A_H2F_A,
       I2C1_SDA_MGPIO0A_H2F_B,
       MDCF,
       MDOENF,
       MDOF,
       MMUART0_CTS_MGPIO19B_H2F_A,
       MMUART0_CTS_MGPIO19B_H2F_B,
       MMUART0_DCD_MGPIO22B_H2F_A,
       MMUART0_DCD_MGPIO22B_H2F_B,
       MMUART0_DSR_MGPIO20B_H2F_A,
       MMUART0_DSR_MGPIO20B_H2F_B,
       MMUART0_DTR_MGPIO18B_H2F_A,
       MMUART0_DTR_MGPIO18B_H2F_B,
       MMUART0_RI_MGPIO21B_H2F_A,
       MMUART0_RI_MGPIO21B_H2F_B,
       MMUART0_RTS_MGPIO17B_H2F_A,
       MMUART0_RTS_MGPIO17B_H2F_B,
       MMUART0_RXD_MGPIO28B_H2F_A,
       MMUART0_RXD_MGPIO28B_H2F_B,
       MMUART0_SCK_MGPIO29B_H2F_A,
       MMUART0_SCK_MGPIO29B_H2F_B,
       MMUART0_TXD_MGPIO27B_H2F_A,
       MMUART0_TXD_MGPIO27B_H2F_B,
       MMUART1_DTR_MGPIO12B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_A,
       MMUART1_RTS_MGPIO11B_H2F_B,
       MMUART1_RXD_MGPIO26B_H2F_A,
       MMUART1_RXD_MGPIO26B_H2F_B,
       MMUART1_SCK_MGPIO25B_H2F_A,
       MMUART1_SCK_MGPIO25B_H2F_B,
       MMUART1_TXD_MGPIO24B_H2F_A,
       MMUART1_TXD_MGPIO24B_H2F_B,
       MPLL_LOCK,
       PER2_FABRIC_PADDR,
       PER2_FABRIC_PENABLE,
       PER2_FABRIC_PSEL,
       PER2_FABRIC_PWDATA,
       PER2_FABRIC_PWRITE,
       RTC_MATCH,
       SLEEPDEEP,
       SLEEPHOLDACK,
       SLEEPING,
       SMBALERT_NO0,
       SMBALERT_NO1,
       SMBSUS_NO0,
       SMBSUS_NO1,
       SPI0_CLK_OUT,
       SPI0_SDI_MGPIO5A_H2F_A,
       SPI0_SDI_MGPIO5A_H2F_B,
       SPI0_SDO_MGPIO6A_H2F_A,
       SPI0_SDO_MGPIO6A_H2F_B,
       SPI0_SS0_MGPIO7A_H2F_A,
       SPI0_SS0_MGPIO7A_H2F_B,
       SPI0_SS1_MGPIO8A_H2F_A,
       SPI0_SS1_MGPIO8A_H2F_B,
       SPI0_SS2_MGPIO9A_H2F_A,
       SPI0_SS2_MGPIO9A_H2F_B,
       SPI0_SS3_MGPIO10A_H2F_A,
       SPI0_SS3_MGPIO10A_H2F_B,
       SPI0_SS4_MGPIO19A_H2F_A,
       SPI0_SS5_MGPIO20A_H2F_A,
       SPI0_SS6_MGPIO21A_H2F_A,
       SPI0_SS7_MGPIO22A_H2F_A,
       SPI1_CLK_OUT,
       SPI1_SDI_MGPIO11A_H2F_A,
       SPI1_SDI_MGPIO11A_H2F_B,
       SPI1_SDO_MGPIO12A_H2F_A,
       SPI1_SDO_MGPIO12A_H2F_B,
       SPI1_SS0_MGPIO13A_H2F_A,
       SPI1_SS0_MGPIO13A_H2F_B,
       SPI1_SS1_MGPIO14A_H2F_A,
       SPI1_SS1_MGPIO14A_H2F_B,
       SPI1_SS2_MGPIO15A_H2F_A,
       SPI1_SS2_MGPIO15A_H2F_B,
       SPI1_SS3_MGPIO16A_H2F_A,
       SPI1_SS3_MGPIO16A_H2F_B,
       SPI1_SS4_MGPIO17A_H2F_A,
       SPI1_SS5_MGPIO18A_H2F_A,
       SPI1_SS6_MGPIO23A_H2F_A,
       SPI1_SS7_MGPIO24A_H2F_A,
       TCGF,
       TRACECLK,
       TRACEDATA,
       TX_CLK,
       TX_ENF,
       TX_ERRF,
       TXCTL_EN_RIF,
       TXD_RIF,
       TXDF,
       TXEV,
       WDOGTIMEOUT,
       F_ARREADY_HREADYOUT1,
       F_AWREADY_HREADYOUT0,
       F_BID,
       F_BRESP_HRESP0,
       F_BVALID,
       F_RDATA_HRDATA01,
       F_RID,
       F_RLAST,
       F_RRESP_HRESP1,
       F_RVALID,
       F_WREADY,
       MDDR_FABRIC_PRDATA,
       MDDR_FABRIC_PREADY,
       MDDR_FABRIC_PSLVERR,
       CAN_RXBUS_F2H_SCP,
       CAN_TX_EBL_F2H_SCP,
       CAN_TXBUS_F2H_SCP,
       COLF,
       CRSF,
       F2_DMAREADY,
       F2H_INTERRUPT,
       F2HCALIB,
       F_DMAREADY,
       F_FM0_ADDR,
       F_FM0_ENABLE,
       F_FM0_MASTLOCK,
       F_FM0_READY,
       F_FM0_SEL,
       F_FM0_SIZE,
       F_FM0_TRANS1,
       F_FM0_WDATA,
       F_FM0_WRITE,
       F_HM0_RDATA,
       F_HM0_READY,
       F_HM0_RESP,
       FAB_AVALID,
       FAB_HOSTDISCON,
       FAB_IDDIG,
       FAB_LINESTATE,
       FAB_M3_RESET_N,
       FAB_PLL_LOCK,
       FAB_RXACTIVE,
       FAB_RXERROR,
       FAB_RXVALID,
       FAB_RXVALIDH,
       FAB_SESSEND,
       FAB_TXREADY,
       FAB_VBUSVALID,
       FAB_VSTATUS,
       FAB_XDATAIN,
       GTX_CLKPF,
       I2C0_BCLK,
       I2C0_SCL_F2H_SCP,
       I2C0_SDA_F2H_SCP,
       I2C1_BCLK,
       I2C1_SCL_F2H_SCP,
       I2C1_SDA_F2H_SCP,
       MDIF,
       MGPIO0A_F2H_GPIN,
       MGPIO10A_F2H_GPIN,
       MGPIO11A_F2H_GPIN,
       MGPIO11B_F2H_GPIN,
       MGPIO12A_F2H_GPIN,
       MGPIO13A_F2H_GPIN,
       MGPIO14A_F2H_GPIN,
       MGPIO15A_F2H_GPIN,
       MGPIO16A_F2H_GPIN,
       MGPIO17B_F2H_GPIN,
       MGPIO18B_F2H_GPIN,
       MGPIO19B_F2H_GPIN,
       MGPIO1A_F2H_GPIN,
       MGPIO20B_F2H_GPIN,
       MGPIO21B_F2H_GPIN,
       MGPIO22B_F2H_GPIN,
       MGPIO24B_F2H_GPIN,
       MGPIO25B_F2H_GPIN,
       MGPIO26B_F2H_GPIN,
       MGPIO27B_F2H_GPIN,
       MGPIO28B_F2H_GPIN,
       MGPIO29B_F2H_GPIN,
       MGPIO2A_F2H_GPIN,
       MGPIO30B_F2H_GPIN,
       MGPIO31B_F2H_GPIN,
       MGPIO3A_F2H_GPIN,
       MGPIO4A_F2H_GPIN,
       MGPIO5A_F2H_GPIN,
       MGPIO6A_F2H_GPIN,
       MGPIO7A_F2H_GPIN,
       MGPIO8A_F2H_GPIN,
       MGPIO9A_F2H_GPIN,
       MMUART0_CTS_F2H_SCP,
       MMUART0_DCD_F2H_SCP,
       MMUART0_DSR_F2H_SCP,
       MMUART0_DTR_F2H_SCP,
       MMUART0_RI_F2H_SCP,
       MMUART0_RTS_F2H_SCP,
       MMUART0_RXD_F2H_SCP,
       MMUART0_SCK_F2H_SCP,
       MMUART0_TXD_F2H_SCP,
       MMUART1_CTS_F2H_SCP,
       MMUART1_DCD_F2H_SCP,
       MMUART1_DSR_F2H_SCP,
       MMUART1_RI_F2H_SCP,
       MMUART1_RTS_F2H_SCP,
       MMUART1_RXD_F2H_SCP,
       MMUART1_SCK_F2H_SCP,
       MMUART1_TXD_F2H_SCP,
       PER2_FABRIC_PRDATA,
       PER2_FABRIC_PREADY,
       PER2_FABRIC_PSLVERR,
       RCGF,
       RX_CLKPF,
       RX_DVF,
       RX_ERRF,
       RX_EV,
       RXDF,
       SLEEPHOLDREQ,
       SMBALERT_NI0,
       SMBALERT_NI1,
       SMBSUS_NI0,
       SMBSUS_NI1,
       SPI0_CLK_IN,
       SPI0_SDI_F2H_SCP,
       SPI0_SDO_F2H_SCP,
       SPI0_SS0_F2H_SCP,
       SPI0_SS1_F2H_SCP,
       SPI0_SS2_F2H_SCP,
       SPI0_SS3_F2H_SCP,
       SPI1_CLK_IN,
       SPI1_SDI_F2H_SCP,
       SPI1_SDO_F2H_SCP,
       SPI1_SS0_F2H_SCP,
       SPI1_SS1_F2H_SCP,
       SPI1_SS2_F2H_SCP,
       SPI1_SS3_F2H_SCP,
       TX_CLKPF,
       USER_MSS_GPIO_RESET_N,
       USER_MSS_RESET_N,
       XCLK_FAB,
       CLK_BASE,
       CLK_MDDR_APB,
       F_ARADDR_HADDR1,
       F_ARBURST_HTRANS1,
       F_ARID_HSEL1,
       F_ARLEN_HBURST1,
       F_ARLOCK_HMASTLOCK1,
       F_ARSIZE_HSIZE1,
       F_ARVALID_HWRITE1,
       F_AWADDR_HADDR0,
       F_AWBURST_HTRANS0,
       F_AWID_HSEL0,
       F_AWLEN_HBURST0,
       F_AWLOCK_HMASTLOCK0,
       F_AWSIZE_HSIZE0,
       F_AWVALID_HWRITE0,
       F_BREADY,
       F_RMW_AXI,
       F_RREADY,
       F_WDATA_HWDATA01,
       F_WID_HREADY01,
       F_WLAST,
       F_WSTRB,
       F_WVALID,
       FPGA_MDDR_ARESET_N,
       MDDR_FABRIC_PADDR,
       MDDR_FABRIC_PENABLE,
       MDDR_FABRIC_PSEL,
       MDDR_FABRIC_PWDATA,
       MDDR_FABRIC_PWRITE,
       PRESET_N,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_IN,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_IN,
       DM_IN,
       DRAM_DQ_IN,
       DRAM_DQS_IN,
       DRAM_FIFO_WE_IN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_IN,
       I2C0_SDA_USBC_DATA0_MGPIO30B_IN,
       I2C1_SCL_USBA_DATA4_MGPIO1A_IN,
       I2C1_SDA_USBA_DATA3_MGPIO0A_IN,
       MGPIO0B_IN,
       MGPIO10B_IN,
       MGPIO1B_IN,
       MGPIO25A_IN,
       MGPIO26A_IN,
       MGPIO27A_IN,
       MGPIO28A_IN,
       MGPIO29A_IN,
       MGPIO2B_IN,
       MGPIO30A_IN,
       MGPIO31A_IN,
       MGPIO3B_IN,
       MGPIO4B_IN,
       MGPIO5B_IN,
       MGPIO6B_IN,
       MGPIO7B_IN,
       MGPIO8B_IN,
       MGPIO9B_IN,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_IN,
       MMUART0_DCD_MGPIO22B_IN,
       MMUART0_DSR_MGPIO20B_IN,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_IN,
       MMUART0_RI_MGPIO21B_IN,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_IN,
       MMUART0_RXD_USBC_STP_MGPIO28B_IN,
       MMUART0_SCK_USBC_NXT_MGPIO29B_IN,
       MMUART0_TXD_USBC_DIR_MGPIO27B_IN,
       MMUART1_CTS_MGPIO13B_IN,
       MMUART1_DCD_MGPIO16B_IN,
       MMUART1_DSR_MGPIO14B_IN,
       MMUART1_DTR_MGPIO12B_IN,
       MMUART1_RI_MGPIO15B_IN,
       MMUART1_RTS_MGPIO11B_IN,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_IN,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_IN,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_IN,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN,
       RGMII_MDC_RMII_MDC_IN,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN,
       RGMII_RX_CLK_IN,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN,
       RGMII_RXD3_USBB_DATA4_IN,
       RGMII_TX_CLK_IN,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_IN,
       RGMII_TXD1_RMII_TXD1_USBB_STP_IN,
       RGMII_TXD2_USBB_DATA5_IN,
       RGMII_TXD3_USBB_DATA6_IN,
       SPI0_SCK_USBA_XCLK_IN,
       SPI0_SDI_USBA_DIR_MGPIO5A_IN,
       SPI0_SDO_USBA_STP_MGPIO6A_IN,
       SPI0_SS0_USBA_NXT_MGPIO7A_IN,
       SPI0_SS1_USBA_DATA5_MGPIO8A_IN,
       SPI0_SS2_USBA_DATA6_MGPIO9A_IN,
       SPI0_SS3_USBA_DATA7_MGPIO10A_IN,
       SPI0_SS4_MGPIO19A_IN,
       SPI0_SS5_MGPIO20A_IN,
       SPI0_SS6_MGPIO21A_IN,
       SPI0_SS7_MGPIO22A_IN,
       SPI1_SCK_IN,
       SPI1_SDI_MGPIO11A_IN,
       SPI1_SDO_MGPIO12A_IN,
       SPI1_SS0_MGPIO13A_IN,
       SPI1_SS1_MGPIO14A_IN,
       SPI1_SS2_MGPIO15A_IN,
       SPI1_SS3_MGPIO16A_IN,
       SPI1_SS4_MGPIO17A_IN,
       SPI1_SS5_MGPIO18A_IN,
       SPI1_SS6_MGPIO23A_IN,
       SPI1_SS7_MGPIO24A_IN,
       USBC_XCLK_IN,
       USBD_DATA0_IN,
       USBD_DATA1_IN,
       USBD_DATA2_IN,
       USBD_DATA3_IN,
       USBD_DATA4_IN,
       USBD_DATA5_IN,
       USBD_DATA6_IN,
       USBD_DATA7_MGPIO23B_IN,
       USBD_DIR_IN,
       USBD_NXT_IN,
       USBD_STP_IN,
       USBD_XCLK_IN,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT,
       DRAM_ADDR,
       DRAM_BA,
       DRAM_CASN,
       DRAM_CKE,
       DRAM_CLK,
       DRAM_CSN,
       DRAM_DM_RDQS_OUT,
       DRAM_DQ_OUT,
       DRAM_DQS_OUT,
       DRAM_FIFO_WE_OUT,
       DRAM_ODT,
       DRAM_RASN,
       DRAM_RSTN,
       DRAM_WEN,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OUT,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OUT,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OUT,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OUT,
       MGPIO0B_OUT,
       MGPIO10B_OUT,
       MGPIO1B_OUT,
       MGPIO25A_OUT,
       MGPIO26A_OUT,
       MGPIO27A_OUT,
       MGPIO28A_OUT,
       MGPIO29A_OUT,
       MGPIO2B_OUT,
       MGPIO30A_OUT,
       MGPIO31A_OUT,
       MGPIO3B_OUT,
       MGPIO4B_OUT,
       MGPIO5B_OUT,
       MGPIO6B_OUT,
       MGPIO7B_OUT,
       MGPIO8B_OUT,
       MGPIO9B_OUT,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT,
       MMUART0_DCD_MGPIO22B_OUT,
       MMUART0_DSR_MGPIO20B_OUT,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT,
       MMUART0_RI_MGPIO21B_OUT,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT,
       MMUART0_RXD_USBC_STP_MGPIO28B_OUT,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OUT,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OUT,
       MMUART1_CTS_MGPIO13B_OUT,
       MMUART1_DCD_MGPIO16B_OUT,
       MMUART1_DSR_MGPIO14B_OUT,
       MMUART1_DTR_MGPIO12B_OUT,
       MMUART1_RI_MGPIO15B_OUT,
       MMUART1_RTS_MGPIO11B_OUT,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT,
       RGMII_MDC_RMII_MDC_OUT,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT,
       RGMII_RX_CLK_OUT,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT,
       RGMII_RXD3_USBB_DATA4_OUT,
       RGMII_TX_CLK_OUT,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OUT,
       RGMII_TXD2_USBB_DATA5_OUT,
       RGMII_TXD3_USBB_DATA6_OUT,
       SPI0_SCK_USBA_XCLK_OUT,
       SPI0_SDI_USBA_DIR_MGPIO5A_OUT,
       SPI0_SDO_USBA_STP_MGPIO6A_OUT,
       SPI0_SS0_USBA_NXT_MGPIO7A_OUT,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OUT,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OUT,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OUT,
       SPI0_SS4_MGPIO19A_OUT,
       SPI0_SS5_MGPIO20A_OUT,
       SPI0_SS6_MGPIO21A_OUT,
       SPI0_SS7_MGPIO22A_OUT,
       SPI1_SCK_OUT,
       SPI1_SDI_MGPIO11A_OUT,
       SPI1_SDO_MGPIO12A_OUT,
       SPI1_SS0_MGPIO13A_OUT,
       SPI1_SS1_MGPIO14A_OUT,
       SPI1_SS2_MGPIO15A_OUT,
       SPI1_SS3_MGPIO16A_OUT,
       SPI1_SS4_MGPIO17A_OUT,
       SPI1_SS5_MGPIO18A_OUT,
       SPI1_SS6_MGPIO23A_OUT,
       SPI1_SS7_MGPIO24A_OUT,
       USBC_XCLK_OUT,
       USBD_DATA0_OUT,
       USBD_DATA1_OUT,
       USBD_DATA2_OUT,
       USBD_DATA3_OUT,
       USBD_DATA4_OUT,
       USBD_DATA5_OUT,
       USBD_DATA6_OUT,
       USBD_DATA7_MGPIO23B_OUT,
       USBD_DIR_OUT,
       USBD_NXT_OUT,
       USBD_STP_OUT,
       USBD_XCLK_OUT,
       CAN_RXBUS_USBA_DATA1_MGPIO3A_OE,
       CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE,
       CAN_TXBUS_USBA_DATA0_MGPIO2A_OE,
       DM_OE,
       DRAM_DQ_OE,
       DRAM_DQS_OE,
       I2C0_SCL_USBC_DATA1_MGPIO31B_OE,
       I2C0_SDA_USBC_DATA0_MGPIO30B_OE,
       I2C1_SCL_USBA_DATA4_MGPIO1A_OE,
       I2C1_SDA_USBA_DATA3_MGPIO0A_OE,
       MGPIO0B_OE,
       MGPIO10B_OE,
       MGPIO1B_OE,
       MGPIO25A_OE,
       MGPIO26A_OE,
       MGPIO27A_OE,
       MGPIO28A_OE,
       MGPIO29A_OE,
       MGPIO2B_OE,
       MGPIO30A_OE,
       MGPIO31A_OE,
       MGPIO3B_OE,
       MGPIO4B_OE,
       MGPIO5B_OE,
       MGPIO6B_OE,
       MGPIO7B_OE,
       MGPIO8B_OE,
       MGPIO9B_OE,
       MMUART0_CTS_USBC_DATA7_MGPIO19B_OE,
       MMUART0_DCD_MGPIO22B_OE,
       MMUART0_DSR_MGPIO20B_OE,
       MMUART0_DTR_USBC_DATA6_MGPIO18B_OE,
       MMUART0_RI_MGPIO21B_OE,
       MMUART0_RTS_USBC_DATA5_MGPIO17B_OE,
       MMUART0_RXD_USBC_STP_MGPIO28B_OE,
       MMUART0_SCK_USBC_NXT_MGPIO29B_OE,
       MMUART0_TXD_USBC_DIR_MGPIO27B_OE,
       MMUART1_CTS_MGPIO13B_OE,
       MMUART1_DCD_MGPIO16B_OE,
       MMUART1_DSR_MGPIO14B_OE,
       MMUART1_DTR_MGPIO12B_OE,
       MMUART1_RI_MGPIO15B_OE,
       MMUART1_RTS_MGPIO11B_OE,
       MMUART1_RXD_USBC_DATA3_MGPIO26B_OE,
       MMUART1_SCK_USBC_DATA4_MGPIO25B_OE,
       MMUART1_TXD_USBC_DATA2_MGPIO24B_OE,
       RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE,
       RGMII_MDC_RMII_MDC_OE,
       RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE,
       RGMII_RX_CLK_OE,
       RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE,
       RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE,
       RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE,
       RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE,
       RGMII_RXD3_USBB_DATA4_OE,
       RGMII_TX_CLK_OE,
       RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE,
       RGMII_TXD0_RMII_TXD0_USBB_DIR_OE,
       RGMII_TXD1_RMII_TXD1_USBB_STP_OE,
       RGMII_TXD2_USBB_DATA5_OE,
       RGMII_TXD3_USBB_DATA6_OE,
       SPI0_SCK_USBA_XCLK_OE,
       SPI0_SDI_USBA_DIR_MGPIO5A_OE,
       SPI0_SDO_USBA_STP_MGPIO6A_OE,
       SPI0_SS0_USBA_NXT_MGPIO7A_OE,
       SPI0_SS1_USBA_DATA5_MGPIO8A_OE,
       SPI0_SS2_USBA_DATA6_MGPIO9A_OE,
       SPI0_SS3_USBA_DATA7_MGPIO10A_OE,
       SPI0_SS4_MGPIO19A_OE,
       SPI0_SS5_MGPIO20A_OE,
       SPI0_SS6_MGPIO21A_OE,
       SPI0_SS7_MGPIO22A_OE,
       SPI1_SCK_OE,
       SPI1_SDI_MGPIO11A_OE,
       SPI1_SDO_MGPIO12A_OE,
       SPI1_SS0_MGPIO13A_OE,
       SPI1_SS1_MGPIO14A_OE,
       SPI1_SS2_MGPIO15A_OE,
       SPI1_SS3_MGPIO16A_OE,
       SPI1_SS4_MGPIO17A_OE,
       SPI1_SS5_MGPIO18A_OE,
       SPI1_SS6_MGPIO23A_OE,
       SPI1_SS7_MGPIO24A_OE,
       USBC_XCLK_OE,
       USBD_DATA0_OE,
       USBD_DATA1_OE,
       USBD_DATA2_OE,
       USBD_DATA3_OE,
       USBD_DATA4_OE,
       USBD_DATA5_OE,
       USBD_DATA6_OE,
       USBD_DATA7_MGPIO23B_OE,
       USBD_DIR_OE,
       USBD_NXT_OE,
       USBD_STP_OE,
       USBD_XCLK_OE
    );
output CAN_RXBUS_MGPIO3A_H2F_A;
output CAN_RXBUS_MGPIO3A_H2F_B;
output CAN_TX_EBL_MGPIO4A_H2F_A;
output CAN_TX_EBL_MGPIO4A_H2F_B;
output CAN_TXBUS_MGPIO2A_H2F_A;
output CAN_TXBUS_MGPIO2A_H2F_B;
output CLK_CONFIG_APB;
output COMMS_INT;
output CONFIG_PRESET_N;
output [7:0] EDAC_ERROR;
output [31:0] F_FM0_RDATA;
output F_FM0_READYOUT;
output F_FM0_RESP;
output [31:0] F_HM0_ADDR;
output F_HM0_ENABLE;
output F_HM0_SEL;
output [1:0] F_HM0_SIZE;
output F_HM0_TRANS1;
output [31:0] F_HM0_WDATA;
output F_HM0_WRITE;
output FAB_CHRGVBUS;
output FAB_DISCHRGVBUS;
output FAB_DMPULLDOWN;
output FAB_DPPULLDOWN;
output FAB_DRVVBUS;
output FAB_IDPULLUP;
output [1:0] FAB_OPMODE;
output FAB_SUSPENDM;
output FAB_TERMSEL;
output FAB_TXVALID;
output [3:0] FAB_VCONTROL;
output FAB_VCONTROLLOADM;
output [1:0] FAB_XCVRSEL;
output [7:0] FAB_XDATAOUT;
output FACC_GLMUX_SEL;
output [1:0] FIC32_0_MASTER;
output [1:0] FIC32_1_MASTER;
output FPGA_RESET_N;
output GTX_CLK;
output [15:0] H2F_INTERRUPT;
output H2F_NMI;
output H2FCALIB;
output I2C0_SCL_MGPIO31B_H2F_A;
output I2C0_SCL_MGPIO31B_H2F_B;
output I2C0_SDA_MGPIO30B_H2F_A;
output I2C0_SDA_MGPIO30B_H2F_B;
output I2C1_SCL_MGPIO1A_H2F_A;
output I2C1_SCL_MGPIO1A_H2F_B;
output I2C1_SDA_MGPIO0A_H2F_A;
output I2C1_SDA_MGPIO0A_H2F_B;
output MDCF;
output MDOENF;
output MDOF;
output MMUART0_CTS_MGPIO19B_H2F_A;
output MMUART0_CTS_MGPIO19B_H2F_B;
output MMUART0_DCD_MGPIO22B_H2F_A;
output MMUART0_DCD_MGPIO22B_H2F_B;
output MMUART0_DSR_MGPIO20B_H2F_A;
output MMUART0_DSR_MGPIO20B_H2F_B;
output MMUART0_DTR_MGPIO18B_H2F_A;
output MMUART0_DTR_MGPIO18B_H2F_B;
output MMUART0_RI_MGPIO21B_H2F_A;
output MMUART0_RI_MGPIO21B_H2F_B;
output MMUART0_RTS_MGPIO17B_H2F_A;
output MMUART0_RTS_MGPIO17B_H2F_B;
output MMUART0_RXD_MGPIO28B_H2F_A;
output MMUART0_RXD_MGPIO28B_H2F_B;
output MMUART0_SCK_MGPIO29B_H2F_A;
output MMUART0_SCK_MGPIO29B_H2F_B;
output MMUART0_TXD_MGPIO27B_H2F_A;
output MMUART0_TXD_MGPIO27B_H2F_B;
output MMUART1_DTR_MGPIO12B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_A;
output MMUART1_RTS_MGPIO11B_H2F_B;
output MMUART1_RXD_MGPIO26B_H2F_A;
output MMUART1_RXD_MGPIO26B_H2F_B;
output MMUART1_SCK_MGPIO25B_H2F_A;
output MMUART1_SCK_MGPIO25B_H2F_B;
output MMUART1_TXD_MGPIO24B_H2F_A;
output MMUART1_TXD_MGPIO24B_H2F_B;
output MPLL_LOCK;
output [15:2] PER2_FABRIC_PADDR;
output PER2_FABRIC_PENABLE;
output PER2_FABRIC_PSEL;
output [31:0] PER2_FABRIC_PWDATA;
output PER2_FABRIC_PWRITE;
output RTC_MATCH;
output SLEEPDEEP;
output SLEEPHOLDACK;
output SLEEPING;
output SMBALERT_NO0;
output SMBALERT_NO1;
output SMBSUS_NO0;
output SMBSUS_NO1;
output SPI0_CLK_OUT;
output SPI0_SDI_MGPIO5A_H2F_A;
output SPI0_SDI_MGPIO5A_H2F_B;
output SPI0_SDO_MGPIO6A_H2F_A;
output SPI0_SDO_MGPIO6A_H2F_B;
output SPI0_SS0_MGPIO7A_H2F_A;
output SPI0_SS0_MGPIO7A_H2F_B;
output SPI0_SS1_MGPIO8A_H2F_A;
output SPI0_SS1_MGPIO8A_H2F_B;
output SPI0_SS2_MGPIO9A_H2F_A;
output SPI0_SS2_MGPIO9A_H2F_B;
output SPI0_SS3_MGPIO10A_H2F_A;
output SPI0_SS3_MGPIO10A_H2F_B;
output SPI0_SS4_MGPIO19A_H2F_A;
output SPI0_SS5_MGPIO20A_H2F_A;
output SPI0_SS6_MGPIO21A_H2F_A;
output SPI0_SS7_MGPIO22A_H2F_A;
output SPI1_CLK_OUT;
output SPI1_SDI_MGPIO11A_H2F_A;
output SPI1_SDI_MGPIO11A_H2F_B;
output SPI1_SDO_MGPIO12A_H2F_A;
output SPI1_SDO_MGPIO12A_H2F_B;
output SPI1_SS0_MGPIO13A_H2F_A;
output SPI1_SS0_MGPIO13A_H2F_B;
output SPI1_SS1_MGPIO14A_H2F_A;
output SPI1_SS1_MGPIO14A_H2F_B;
output SPI1_SS2_MGPIO15A_H2F_A;
output SPI1_SS2_MGPIO15A_H2F_B;
output SPI1_SS3_MGPIO16A_H2F_A;
output SPI1_SS3_MGPIO16A_H2F_B;
output SPI1_SS4_MGPIO17A_H2F_A;
output SPI1_SS5_MGPIO18A_H2F_A;
output SPI1_SS6_MGPIO23A_H2F_A;
output SPI1_SS7_MGPIO24A_H2F_A;
output [9:0] TCGF;
output TRACECLK;
output [3:0] TRACEDATA;
output TX_CLK;
output TX_ENF;
output TX_ERRF;
output TXCTL_EN_RIF;
output [3:0] TXD_RIF;
output [7:0] TXDF;
output TXEV;
output WDOGTIMEOUT;
output F_ARREADY_HREADYOUT1;
output F_AWREADY_HREADYOUT0;
output [3:0] F_BID;
output [1:0] F_BRESP_HRESP0;
output F_BVALID;
output [63:0] F_RDATA_HRDATA01;
output [3:0] F_RID;
output F_RLAST;
output [1:0] F_RRESP_HRESP1;
output F_RVALID;
output F_WREADY;
output [15:0] MDDR_FABRIC_PRDATA;
output MDDR_FABRIC_PREADY;
output MDDR_FABRIC_PSLVERR;
input  CAN_RXBUS_F2H_SCP;
input  CAN_TX_EBL_F2H_SCP;
input  CAN_TXBUS_F2H_SCP;
input  COLF;
input  CRSF;
input  [1:0] F2_DMAREADY;
input  [15:0] F2H_INTERRUPT;
input  F2HCALIB;
input  [1:0] F_DMAREADY;
input  [31:0] F_FM0_ADDR;
input  F_FM0_ENABLE;
input  F_FM0_MASTLOCK;
input  F_FM0_READY;
input  F_FM0_SEL;
input  [1:0] F_FM0_SIZE;
input  F_FM0_TRANS1;
input  [31:0] F_FM0_WDATA;
input  F_FM0_WRITE;
input  [31:0] F_HM0_RDATA;
input  F_HM0_READY;
input  F_HM0_RESP;
input  FAB_AVALID;
input  FAB_HOSTDISCON;
input  FAB_IDDIG;
input  [1:0] FAB_LINESTATE;
input  FAB_M3_RESET_N;
input  FAB_PLL_LOCK;
input  FAB_RXACTIVE;
input  FAB_RXERROR;
input  FAB_RXVALID;
input  FAB_RXVALIDH;
input  FAB_SESSEND;
input  FAB_TXREADY;
input  FAB_VBUSVALID;
input  [7:0] FAB_VSTATUS;
input  [7:0] FAB_XDATAIN;
input  GTX_CLKPF;
input  I2C0_BCLK;
input  I2C0_SCL_F2H_SCP;
input  I2C0_SDA_F2H_SCP;
input  I2C1_BCLK;
input  I2C1_SCL_F2H_SCP;
input  I2C1_SDA_F2H_SCP;
input  MDIF;
input  MGPIO0A_F2H_GPIN;
input  MGPIO10A_F2H_GPIN;
input  MGPIO11A_F2H_GPIN;
input  MGPIO11B_F2H_GPIN;
input  MGPIO12A_F2H_GPIN;
input  MGPIO13A_F2H_GPIN;
input  MGPIO14A_F2H_GPIN;
input  MGPIO15A_F2H_GPIN;
input  MGPIO16A_F2H_GPIN;
input  MGPIO17B_F2H_GPIN;
input  MGPIO18B_F2H_GPIN;
input  MGPIO19B_F2H_GPIN;
input  MGPIO1A_F2H_GPIN;
input  MGPIO20B_F2H_GPIN;
input  MGPIO21B_F2H_GPIN;
input  MGPIO22B_F2H_GPIN;
input  MGPIO24B_F2H_GPIN;
input  MGPIO25B_F2H_GPIN;
input  MGPIO26B_F2H_GPIN;
input  MGPIO27B_F2H_GPIN;
input  MGPIO28B_F2H_GPIN;
input  MGPIO29B_F2H_GPIN;
input  MGPIO2A_F2H_GPIN;
input  MGPIO30B_F2H_GPIN;
input  MGPIO31B_F2H_GPIN;
input  MGPIO3A_F2H_GPIN;
input  MGPIO4A_F2H_GPIN;
input  MGPIO5A_F2H_GPIN;
input  MGPIO6A_F2H_GPIN;
input  MGPIO7A_F2H_GPIN;
input  MGPIO8A_F2H_GPIN;
input  MGPIO9A_F2H_GPIN;
input  MMUART0_CTS_F2H_SCP;
input  MMUART0_DCD_F2H_SCP;
input  MMUART0_DSR_F2H_SCP;
input  MMUART0_DTR_F2H_SCP;
input  MMUART0_RI_F2H_SCP;
input  MMUART0_RTS_F2H_SCP;
input  MMUART0_RXD_F2H_SCP;
input  MMUART0_SCK_F2H_SCP;
input  MMUART0_TXD_F2H_SCP;
input  MMUART1_CTS_F2H_SCP;
input  MMUART1_DCD_F2H_SCP;
input  MMUART1_DSR_F2H_SCP;
input  MMUART1_RI_F2H_SCP;
input  MMUART1_RTS_F2H_SCP;
input  MMUART1_RXD_F2H_SCP;
input  MMUART1_SCK_F2H_SCP;
input  MMUART1_TXD_F2H_SCP;
input  [31:0] PER2_FABRIC_PRDATA;
input  PER2_FABRIC_PREADY;
input  PER2_FABRIC_PSLVERR;
input  [9:0] RCGF;
input  RX_CLKPF;
input  RX_DVF;
input  RX_ERRF;
input  RX_EV;
input  [7:0] RXDF;
input  SLEEPHOLDREQ;
input  SMBALERT_NI0;
input  SMBALERT_NI1;
input  SMBSUS_NI0;
input  SMBSUS_NI1;
input  SPI0_CLK_IN;
input  SPI0_SDI_F2H_SCP;
input  SPI0_SDO_F2H_SCP;
input  SPI0_SS0_F2H_SCP;
input  SPI0_SS1_F2H_SCP;
input  SPI0_SS2_F2H_SCP;
input  SPI0_SS3_F2H_SCP;
input  SPI1_CLK_IN;
input  SPI1_SDI_F2H_SCP;
input  SPI1_SDO_F2H_SCP;
input  SPI1_SS0_F2H_SCP;
input  SPI1_SS1_F2H_SCP;
input  SPI1_SS2_F2H_SCP;
input  SPI1_SS3_F2H_SCP;
input  TX_CLKPF;
input  USER_MSS_GPIO_RESET_N;
input  USER_MSS_RESET_N;
input  XCLK_FAB;
input  CLK_BASE;
input  CLK_MDDR_APB;
input  [31:0] F_ARADDR_HADDR1;
input  [1:0] F_ARBURST_HTRANS1;
input  [3:0] F_ARID_HSEL1;
input  [3:0] F_ARLEN_HBURST1;
input  [1:0] F_ARLOCK_HMASTLOCK1;
input  [1:0] F_ARSIZE_HSIZE1;
input  F_ARVALID_HWRITE1;
input  [31:0] F_AWADDR_HADDR0;
input  [1:0] F_AWBURST_HTRANS0;
input  [3:0] F_AWID_HSEL0;
input  [3:0] F_AWLEN_HBURST0;
input  [1:0] F_AWLOCK_HMASTLOCK0;
input  [1:0] F_AWSIZE_HSIZE0;
input  F_AWVALID_HWRITE0;
input  F_BREADY;
input  F_RMW_AXI;
input  F_RREADY;
input  [63:0] F_WDATA_HWDATA01;
input  [3:0] F_WID_HREADY01;
input  F_WLAST;
input  [7:0] F_WSTRB;
input  F_WVALID;
input  FPGA_MDDR_ARESET_N;
input  [10:2] MDDR_FABRIC_PADDR;
input  MDDR_FABRIC_PENABLE;
input  MDDR_FABRIC_PSEL;
input  [15:0] MDDR_FABRIC_PWDATA;
input  MDDR_FABRIC_PWRITE;
input  PRESET_N;
input  CAN_RXBUS_USBA_DATA1_MGPIO3A_IN;
input  CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN;
input  CAN_TXBUS_USBA_DATA0_MGPIO2A_IN;
input  [2:0] DM_IN;
input  [17:0] DRAM_DQ_IN;
input  [2:0] DRAM_DQS_IN;
input  [1:0] DRAM_FIFO_WE_IN;
input  I2C0_SCL_USBC_DATA1_MGPIO31B_IN;
input  I2C0_SDA_USBC_DATA0_MGPIO30B_IN;
input  I2C1_SCL_USBA_DATA4_MGPIO1A_IN;
input  I2C1_SDA_USBA_DATA3_MGPIO0A_IN;
input  MGPIO0B_IN;
input  MGPIO10B_IN;
input  MGPIO1B_IN;
input  MGPIO25A_IN;
input  MGPIO26A_IN;
input  MGPIO27A_IN;
input  MGPIO28A_IN;
input  MGPIO29A_IN;
input  MGPIO2B_IN;
input  MGPIO30A_IN;
input  MGPIO31A_IN;
input  MGPIO3B_IN;
input  MGPIO4B_IN;
input  MGPIO5B_IN;
input  MGPIO6B_IN;
input  MGPIO7B_IN;
input  MGPIO8B_IN;
input  MGPIO9B_IN;
input  MMUART0_CTS_USBC_DATA7_MGPIO19B_IN;
input  MMUART0_DCD_MGPIO22B_IN;
input  MMUART0_DSR_MGPIO20B_IN;
input  MMUART0_DTR_USBC_DATA6_MGPIO18B_IN;
input  MMUART0_RI_MGPIO21B_IN;
input  MMUART0_RTS_USBC_DATA5_MGPIO17B_IN;
input  MMUART0_RXD_USBC_STP_MGPIO28B_IN;
input  MMUART0_SCK_USBC_NXT_MGPIO29B_IN;
input  MMUART0_TXD_USBC_DIR_MGPIO27B_IN;
input  MMUART1_CTS_MGPIO13B_IN;
input  MMUART1_DCD_MGPIO16B_IN;
input  MMUART1_DSR_MGPIO14B_IN;
input  MMUART1_DTR_MGPIO12B_IN;
input  MMUART1_RI_MGPIO15B_IN;
input  MMUART1_RTS_MGPIO11B_IN;
input  MMUART1_RXD_USBC_DATA3_MGPIO26B_IN;
input  MMUART1_SCK_USBC_DATA4_MGPIO25B_IN;
input  MMUART1_TXD_USBC_DATA2_MGPIO24B_IN;
input  RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN;
input  RGMII_MDC_RMII_MDC_IN;
input  RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN;
input  RGMII_RX_CLK_IN;
input  RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN;
input  RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN;
input  RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN;
input  RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN;
input  RGMII_RXD3_USBB_DATA4_IN;
input  RGMII_TX_CLK_IN;
input  RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN;
input  RGMII_TXD0_RMII_TXD0_USBB_DIR_IN;
input  RGMII_TXD1_RMII_TXD1_USBB_STP_IN;
input  RGMII_TXD2_USBB_DATA5_IN;
input  RGMII_TXD3_USBB_DATA6_IN;
input  SPI0_SCK_USBA_XCLK_IN;
input  SPI0_SDI_USBA_DIR_MGPIO5A_IN;
input  SPI0_SDO_USBA_STP_MGPIO6A_IN;
input  SPI0_SS0_USBA_NXT_MGPIO7A_IN;
input  SPI0_SS1_USBA_DATA5_MGPIO8A_IN;
input  SPI0_SS2_USBA_DATA6_MGPIO9A_IN;
input  SPI0_SS3_USBA_DATA7_MGPIO10A_IN;
input  SPI0_SS4_MGPIO19A_IN;
input  SPI0_SS5_MGPIO20A_IN;
input  SPI0_SS6_MGPIO21A_IN;
input  SPI0_SS7_MGPIO22A_IN;
input  SPI1_SCK_IN;
input  SPI1_SDI_MGPIO11A_IN;
input  SPI1_SDO_MGPIO12A_IN;
input  SPI1_SS0_MGPIO13A_IN;
input  SPI1_SS1_MGPIO14A_IN;
input  SPI1_SS2_MGPIO15A_IN;
input  SPI1_SS3_MGPIO16A_IN;
input  SPI1_SS4_MGPIO17A_IN;
input  SPI1_SS5_MGPIO18A_IN;
input  SPI1_SS6_MGPIO23A_IN;
input  SPI1_SS7_MGPIO24A_IN;
input  USBC_XCLK_IN;
input  USBD_DATA0_IN;
input  USBD_DATA1_IN;
input  USBD_DATA2_IN;
input  USBD_DATA3_IN;
input  USBD_DATA4_IN;
input  USBD_DATA5_IN;
input  USBD_DATA6_IN;
input  USBD_DATA7_MGPIO23B_IN;
input  USBD_DIR_IN;
input  USBD_NXT_IN;
input  USBD_STP_IN;
input  USBD_XCLK_IN;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT;
output [15:0] DRAM_ADDR;
output [2:0] DRAM_BA;
output DRAM_CASN;
output DRAM_CKE;
output DRAM_CLK;
output DRAM_CSN;
output [2:0] DRAM_DM_RDQS_OUT;
output [17:0] DRAM_DQ_OUT;
output [2:0] DRAM_DQS_OUT;
output [1:0] DRAM_FIFO_WE_OUT;
output DRAM_ODT;
output DRAM_RASN;
output DRAM_RSTN;
output DRAM_WEN;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OUT;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OUT;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OUT;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OUT;
output MGPIO0B_OUT;
output MGPIO10B_OUT;
output MGPIO1B_OUT;
output MGPIO25A_OUT;
output MGPIO26A_OUT;
output MGPIO27A_OUT;
output MGPIO28A_OUT;
output MGPIO29A_OUT;
output MGPIO2B_OUT;
output MGPIO30A_OUT;
output MGPIO31A_OUT;
output MGPIO3B_OUT;
output MGPIO4B_OUT;
output MGPIO5B_OUT;
output MGPIO6B_OUT;
output MGPIO7B_OUT;
output MGPIO8B_OUT;
output MGPIO9B_OUT;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT;
output MMUART0_DCD_MGPIO22B_OUT;
output MMUART0_DSR_MGPIO20B_OUT;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT;
output MMUART0_RI_MGPIO21B_OUT;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT;
output MMUART0_RXD_USBC_STP_MGPIO28B_OUT;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OUT;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OUT;
output MMUART1_CTS_MGPIO13B_OUT;
output MMUART1_DCD_MGPIO16B_OUT;
output MMUART1_DSR_MGPIO14B_OUT;
output MMUART1_DTR_MGPIO12B_OUT;
output MMUART1_RI_MGPIO15B_OUT;
output MMUART1_RTS_MGPIO11B_OUT;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT;
output RGMII_MDC_RMII_MDC_OUT;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT;
output RGMII_RX_CLK_OUT;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT;
output RGMII_RXD3_USBB_DATA4_OUT;
output RGMII_TX_CLK_OUT;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OUT;
output RGMII_TXD2_USBB_DATA5_OUT;
output RGMII_TXD3_USBB_DATA6_OUT;
output SPI0_SCK_USBA_XCLK_OUT;
output SPI0_SDI_USBA_DIR_MGPIO5A_OUT;
output SPI0_SDO_USBA_STP_MGPIO6A_OUT;
output SPI0_SS0_USBA_NXT_MGPIO7A_OUT;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OUT;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OUT;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OUT;
output SPI0_SS4_MGPIO19A_OUT;
output SPI0_SS5_MGPIO20A_OUT;
output SPI0_SS6_MGPIO21A_OUT;
output SPI0_SS7_MGPIO22A_OUT;
output SPI1_SCK_OUT;
output SPI1_SDI_MGPIO11A_OUT;
output SPI1_SDO_MGPIO12A_OUT;
output SPI1_SS0_MGPIO13A_OUT;
output SPI1_SS1_MGPIO14A_OUT;
output SPI1_SS2_MGPIO15A_OUT;
output SPI1_SS3_MGPIO16A_OUT;
output SPI1_SS4_MGPIO17A_OUT;
output SPI1_SS5_MGPIO18A_OUT;
output SPI1_SS6_MGPIO23A_OUT;
output SPI1_SS7_MGPIO24A_OUT;
output USBC_XCLK_OUT;
output USBD_DATA0_OUT;
output USBD_DATA1_OUT;
output USBD_DATA2_OUT;
output USBD_DATA3_OUT;
output USBD_DATA4_OUT;
output USBD_DATA5_OUT;
output USBD_DATA6_OUT;
output USBD_DATA7_MGPIO23B_OUT;
output USBD_DIR_OUT;
output USBD_NXT_OUT;
output USBD_STP_OUT;
output USBD_XCLK_OUT;
output CAN_RXBUS_USBA_DATA1_MGPIO3A_OE;
output CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE;
output CAN_TXBUS_USBA_DATA0_MGPIO2A_OE;
output [2:0] DM_OE;
output [17:0] DRAM_DQ_OE;
output [2:0] DRAM_DQS_OE;
output I2C0_SCL_USBC_DATA1_MGPIO31B_OE;
output I2C0_SDA_USBC_DATA0_MGPIO30B_OE;
output I2C1_SCL_USBA_DATA4_MGPIO1A_OE;
output I2C1_SDA_USBA_DATA3_MGPIO0A_OE;
output MGPIO0B_OE;
output MGPIO10B_OE;
output MGPIO1B_OE;
output MGPIO25A_OE;
output MGPIO26A_OE;
output MGPIO27A_OE;
output MGPIO28A_OE;
output MGPIO29A_OE;
output MGPIO2B_OE;
output MGPIO30A_OE;
output MGPIO31A_OE;
output MGPIO3B_OE;
output MGPIO4B_OE;
output MGPIO5B_OE;
output MGPIO6B_OE;
output MGPIO7B_OE;
output MGPIO8B_OE;
output MGPIO9B_OE;
output MMUART0_CTS_USBC_DATA7_MGPIO19B_OE;
output MMUART0_DCD_MGPIO22B_OE;
output MMUART0_DSR_MGPIO20B_OE;
output MMUART0_DTR_USBC_DATA6_MGPIO18B_OE;
output MMUART0_RI_MGPIO21B_OE;
output MMUART0_RTS_USBC_DATA5_MGPIO17B_OE;
output MMUART0_RXD_USBC_STP_MGPIO28B_OE;
output MMUART0_SCK_USBC_NXT_MGPIO29B_OE;
output MMUART0_TXD_USBC_DIR_MGPIO27B_OE;
output MMUART1_CTS_MGPIO13B_OE;
output MMUART1_DCD_MGPIO16B_OE;
output MMUART1_DSR_MGPIO14B_OE;
output MMUART1_DTR_MGPIO12B_OE;
output MMUART1_RI_MGPIO15B_OE;
output MMUART1_RTS_MGPIO11B_OE;
output MMUART1_RXD_USBC_DATA3_MGPIO26B_OE;
output MMUART1_SCK_USBC_DATA4_MGPIO25B_OE;
output MMUART1_TXD_USBC_DATA2_MGPIO24B_OE;
output RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE;
output RGMII_MDC_RMII_MDC_OE;
output RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE;
output RGMII_RX_CLK_OE;
output RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE;
output RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE;
output RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE;
output RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE;
output RGMII_RXD3_USBB_DATA4_OE;
output RGMII_TX_CLK_OE;
output RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE;
output RGMII_TXD0_RMII_TXD0_USBB_DIR_OE;
output RGMII_TXD1_RMII_TXD1_USBB_STP_OE;
output RGMII_TXD2_USBB_DATA5_OE;
output RGMII_TXD3_USBB_DATA6_OE;
output SPI0_SCK_USBA_XCLK_OE;
output SPI0_SDI_USBA_DIR_MGPIO5A_OE;
output SPI0_SDO_USBA_STP_MGPIO6A_OE;
output SPI0_SS0_USBA_NXT_MGPIO7A_OE;
output SPI0_SS1_USBA_DATA5_MGPIO8A_OE;
output SPI0_SS2_USBA_DATA6_MGPIO9A_OE;
output SPI0_SS3_USBA_DATA7_MGPIO10A_OE;
output SPI0_SS4_MGPIO19A_OE;
output SPI0_SS5_MGPIO20A_OE;
output SPI0_SS6_MGPIO21A_OE;
output SPI0_SS7_MGPIO22A_OE;
output SPI1_SCK_OE;
output SPI1_SDI_MGPIO11A_OE;
output SPI1_SDO_MGPIO12A_OE;
output SPI1_SS0_MGPIO13A_OE;
output SPI1_SS1_MGPIO14A_OE;
output SPI1_SS2_MGPIO15A_OE;
output SPI1_SS3_MGPIO16A_OE;
output SPI1_SS4_MGPIO17A_OE;
output SPI1_SS5_MGPIO18A_OE;
output SPI1_SS6_MGPIO23A_OE;
output SPI1_SS7_MGPIO24A_OE;
output USBC_XCLK_OE;
output USBD_DATA0_OE;
output USBD_DATA1_OE;
output USBD_DATA2_OE;
output USBD_DATA3_OE;
output USBD_DATA4_OE;
output USBD_DATA5_OE;
output USBD_DATA6_OE;
output USBD_DATA7_MGPIO23B_OE;
output USBD_DIR_OE;
output USBD_NXT_OE;
output USBD_STP_OE;
output USBD_XCLK_OE;

    parameter INIT = 'h0 ;
    parameter ACT_UBITS = 'hFFFFFFFFFFFFFF ;
    parameter MEMORYFILE = "" ;
    parameter RTC_MAIN_XTL_FREQ = 0.0 ;
    parameter RTC_MAIN_XTL_MODE = "1" ;
    parameter DDR_CLK_FREQ = 0.0 ;
    
endmodule


module Ram_intferface(
       TPSRAM_0_RD,
       Ram_intferface_0_o_TPSRAM_WD,
       Ram_intferface_0_o_TPSRAM_RADDR_sv,
       Ram_intferface_0_o_TPSRAM_WADDR_sv,
       Ram_intferface_0_o_TPSRAM_REN,
       Ram_intferface_0_o_TPSRAM_WEN,
       Ram_intferface_0_o_reset_n,
       demo_0_FAB_CCC_GL0,
       demo_0_POWER_ON_RESET_N
    );
input  [7:0] TPSRAM_0_RD;
output [7:0] Ram_intferface_0_o_TPSRAM_WD;
output [5:0] Ram_intferface_0_o_TPSRAM_RADDR_sv;
output [5:0] Ram_intferface_0_o_TPSRAM_WADDR_sv;
output Ram_intferface_0_o_TPSRAM_REN;
output Ram_intferface_0_o_TPSRAM_WEN;
output Ram_intferface_0_o_reset_n;
input  demo_0_FAB_CCC_GL0;
input  demo_0_POWER_ON_RESET_N;

    wire VCC_net_1, \o_TPSRAM_WD_3[5]_net_1 , N_103_i, GND_net_1, 
        \o_TPSRAM_WD_3[6]_net_1 , \o_TPSRAM_WD_3[7]_net_1 , 
        \o_TPSRAM_WADDR_sv_3[0]_net_1 , \o_TPSRAM_WADDR_sv_3[1]_net_1 , 
        \o_TPSRAM_WADDR_sv_3[2]_net_1 , \o_TPSRAM_WADDR_sv_3[3]_net_1 , 
        \o_TPSRAM_WADDR_sv_3[4]_net_1 , \o_TPSRAM_WADDR_sv_3[5]_net_1 , 
        \next_addr[2]_net_1 , \next_addr_6[2]_net_1 , 
        un1_state_tpsram_access_2_0_a3_net_1, \next_addr[3]_net_1 , 
        \next_addr_6[3]_net_1 , \next_addr[4]_net_1 , 
        \next_addr_6[4]_net_1 , \next_addr[5]_net_1 , 
        \next_addr_6[5]_net_1 , \o_TPSRAM_RADDR_sv_6[0]_net_1 , 
        un1_state_tpsram_access_9_0_net_1, 
        \o_TPSRAM_RADDR_sv_6[1]_net_1 , \o_TPSRAM_RADDR_sv_6[2]_net_1 , 
        \o_TPSRAM_RADDR_sv_6[3]_net_1 , \o_TPSRAM_RADDR_sv_6[4]_net_1 , 
        \o_TPSRAM_RADDR_sv_6[5]_net_1 , \o_TPSRAM_WD_3[0]_net_1 , 
        \o_TPSRAM_WD_3[1]_net_1 , \o_TPSRAM_WD_3[2]_net_1 , 
        \o_TPSRAM_WD_3[3]_net_1 , \o_TPSRAM_WD_3[4]_net_1 , 
        \next_addr[0]_net_1 , \next_addr_6[0]_net_1 , 
        \next_addr[1]_net_1 , \next_addr_6[1]_net_1 , 
        \state_tpsram_access[0]_net_1 , un1_state_tpsram_access_7_i, 
        N_90_i, \un1_state_tpsram_access_4[0] , un15_0_net_1, 
        \state_tpsram_access[1]_net_1 , 
        \state_tpsram_access_ns[1]_net_1 , 
        \state_tpsram_access[2]_net_1 , N_76_i, 
        \state_tpsram_access[3]_net_1 , \state_tpsram_access_ns[3] , 
        \state_tpsram_access[4]_net_1 , 
        \state_tpsram_access_ns[4]_net_1 , 
        \state_tpsram_access[5]_net_1 , 
        \state_tpsram_access_ns_a3[5]_net_1 , \next_data[0]_net_1 , 
        \next_data_s[0] , next_datae, \next_data[1]_net_1 , 
        \next_data_s[1] , \next_data[2]_net_1 , \next_data_s[2] , 
        \next_data[3]_net_1 , \next_data_s[3] , \next_data[4]_net_1 , 
        \next_data_s[4] , \next_data[5]_net_1 , \next_data_s[5] , 
        \next_data[6]_net_1 , \next_data_s[6] , \next_data[7]_net_1 , 
        \next_data_s[7]_net_1 , \expected_data[0]_net_1 , 
        \expected_data_s[0] , expected_datae, \expected_data[1]_net_1 , 
        \expected_data_s[1] , \expected_data[2]_net_1 , 
        \expected_data_s[2] , \expected_data[3]_net_1 , 
        \expected_data_s[3] , \expected_data[4]_net_1 , 
        \expected_data_s[4] , \expected_data[5]_net_1 , 
        \expected_data_s[5] , \expected_data[6]_net_1 , 
        \expected_data_s[6] , \expected_data[7]_net_1 , 
        \expected_data_s[7] , \counter[0]_net_1 , \counter_s[0] , 
        countere, \counter[1]_net_1 , \counter_s[1] , 
        \counter[2]_net_1 , \counter_s[2] , \counter[3]_net_1 , 
        \counter_s[3] , \counter[4]_net_1 , \counter_s[4] , 
        \counter[5]_net_1 , \counter_s[5] , \counter[6]_net_1 , 
        \counter_s[6] , \counter[7]_net_1 , \counter_s[7] , 
        \counter[8]_net_1 , \counter_s[8] , \counter[9]_net_1 , 
        \counter_s[9] , \counter[10]_net_1 , \counter_s[10] , 
        \counter[11]_net_1 , \counter_s[11] , \counter[12]_net_1 , 
        \counter_s[12] , \counter[13]_net_1 , \counter_s[13] , 
        \counter[14]_net_1 , \counter_s[14] , \counter[15]_net_1 , 
        \counter_s[15]_net_1 , next_data_cry_cy, 
        \next_data_cry[0]_net_1 , \next_data_cry[1]_net_1 , 
        \next_data_cry[2]_net_1 , \next_data_cry[3]_net_1 , 
        \next_data_cry[4]_net_1 , \next_data_cry[5]_net_1 , 
        \next_data_cry[6]_net_1 , expected_data_cry_cy, 
        o_TPSRAM_WEN8_RNITP5V_Y, o_TPSRAM_WEN8_net_1, 
        \expected_data_cry[0] , \expected_data_cry[1] , 
        \expected_data_cry[2] , \expected_data_cry[3] , 
        \expected_data_cry[4] , \expected_data_cry[5] , 
        \expected_data_cry[6] , counter_cry_cy, \counter_cry[0]_net_1 , 
        \counter_cry[1]_net_1 , \counter_cry[2]_net_1 , 
        \counter_cry[3]_net_1 , \counter_cry[4]_net_1 , 
        \counter_cry[5]_net_1 , \counter_cry[6]_net_1 , 
        \counter_cry[7]_net_1 , \counter_cry[8]_net_1 , 
        \counter_cry[9]_net_1 , \counter_cry[10]_net_1 , 
        \counter_cry[11]_net_1 , \counter_cry[12]_net_1 , 
        \counter_cry[13]_net_1 , \counter_cry[14]_net_1 , 
        o_TPSRAM_WEN8_1_net_1, o_TPSRAM_WEN8_2_net_1, 
        un1_i_TPSRAM_RD_sv_NE_3_net_1, un1_i_TPSRAM_RD_sv_NE_2_net_1, 
        un1_i_TPSRAM_RD_sv_NE_1_net_1, un1_i_TPSRAM_RD_sv_NE_0_net_1, 
        un2_flag_1ms_11_net_1, un2_flag_1ms_10_net_1, 
        un2_flag_1ms_9_net_1, un2_flag_1ms_8_net_1, un6_next_addr_c4, 
        un1_i_TPSRAM_RD_sv_NE_net_1, N_46, un1_state_tpsram_access_10;
    
    SLE \expected_data[0]  (.D(\expected_data_s[0] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[0]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[3]  (.A(VCC_net_1), .B(
        \counter[3]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[2]_net_1 ), .S(\counter_s[3] ), 
        .Y(), .FCO(\counter_cry[3]_net_1 ));
    SLE \o_TPSRAM_WADDR_sv[1]  (.D(\o_TPSRAM_WADDR_sv_3[1]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[1]));
    CFG3 #( .INIT(8'hCA) )  o_reset_n_RNO (.A(
        \state_tpsram_access[0]_net_1 ), .B(
        un1_i_TPSRAM_RD_sv_NE_net_1), .C(
        \state_tpsram_access[4]_net_1 ), .Y(
        un1_state_tpsram_access_7_i));
    SLE \o_TPSRAM_WD[0]  (.D(\o_TPSRAM_WD_3[0]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[0]));
    CFG4 #( .INIT(16'hF1F0) )  \state_tpsram_access_ns[4]  (.A(
        o_TPSRAM_WEN8_net_1), .B(un1_i_TPSRAM_RD_sv_NE_net_1), .C(
        \state_tpsram_access[3]_net_1 ), .D(
        \state_tpsram_access[4]_net_1 ), .Y(
        \state_tpsram_access_ns[4]_net_1 ));
    SLE \state_tpsram_access[2]  (.D(N_76_i), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(VCC_net_1), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[2]_net_1 ));
    SLE \next_addr[0]  (.D(\next_addr_6[0]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[0]_net_1 ));
    SLE \o_TPSRAM_WD[4]  (.D(\o_TPSRAM_WD_3[4]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[4]));
    SLE \next_data[4]  (.D(\next_data_s[4] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[4]_net_1 ));
    CFG4 #( .INIT(16'hCFEF) )  un1_state_tpsram_access_9_0 (.A(
        \state_tpsram_access[4]_net_1 ), .B(
        \state_tpsram_access[3]_net_1 ), .C(o_TPSRAM_WEN8_RNITP5V_Y), 
        .D(o_TPSRAM_WEN8_net_1), .Y(un1_state_tpsram_access_9_0_net_1));
    SLE \counter[11]  (.D(\counter_s[11] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[11]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[3]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[3]_net_1 ), .Y(
        \o_TPSRAM_WD_3[3]_net_1 ));
    SLE \o_TPSRAM_RADDR_sv[5]  (.D(\o_TPSRAM_RADDR_sv_6[5]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[5]));
    SLE \o_TPSRAM_WADDR_sv[2]  (.D(\o_TPSRAM_WADDR_sv_3[2]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[2]));
    SLE \expected_data[1]  (.D(\expected_data_s[1] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[1]_net_1 ));
    SLE \o_TPSRAM_WADDR_sv[3]  (.D(\o_TPSRAM_WADDR_sv_3[3]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[3]));
    CFG4 #( .INIT(16'h0001) )  un2_flag_1ms_9 (.A(\counter[9]_net_1 ), 
        .B(\counter[6]_net_1 ), .C(\counter[4]_net_1 ), .D(
        \counter[2]_net_1 ), .Y(un2_flag_1ms_9_net_1));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[1]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[1]_net_1 ), .Y(
        \o_TPSRAM_WD_3[1]_net_1 ));
    SLE \o_TPSRAM_WD[6]  (.D(\o_TPSRAM_WD_3[6]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[6]));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[6]  (.A(VCC_net_1), .B(
        \next_data[6]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[5]_net_1 ), .S(
        \next_data_s[6] ), .Y(), .FCO(\next_data_cry[6]_net_1 ));
    CFG4 #( .INIT(16'h1000) )  o_TPSRAM_WEN8 (.A(\next_addr[2]_net_1 ), 
        .B(\next_addr[5]_net_1 ), .C(o_TPSRAM_WEN8_2_net_1), .D(
        o_TPSRAM_WEN8_1_net_1), .Y(o_TPSRAM_WEN8_net_1));
    SLE \next_addr[4]  (.D(\next_addr_6[4]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[4]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNIMPL08[5]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[5]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[4] ), .S(\expected_data_s[5] ), .Y(), .FCO(
        \expected_data_cry[5] ));
    CFG3 #( .INIT(8'hBA) )  \state_tpsram_access_ns[1]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(N_46), .C(
        \state_tpsram_access[1]_net_1 ), .Y(
        \state_tpsram_access_ns[1]_net_1 ));
    SLE \counter[6]  (.D(\counter_s[6] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[6]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNIC0BA3[1]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[1]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[0] ), .S(\expected_data_s[1] ), .Y(), .FCO(
        \expected_data_cry[1] ));
    SLE \next_data[5]  (.D(\next_data_s[5] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[5]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  un2_flag_1ms_8 (.A(\counter[15]_net_1 ), 
        .B(\counter[12]_net_1 ), .C(\counter[11]_net_1 ), .D(
        \counter[10]_net_1 ), .Y(un2_flag_1ms_8_net_1));
    SLE \expected_data[4]  (.D(\expected_data_s[4] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[4]_net_1 ));
    SLE \o_TPSRAM_WD[7]  (.D(\o_TPSRAM_WD_3[7]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[7]));
    SLE \counter[3]  (.D(\counter_s[3] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[3]_net_1 ));
    SLE \counter[2]  (.D(\counter_s[2] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[2]_net_1 ));
    CFG3 #( .INIT(8'h48) )  \o_TPSRAM_RADDR_sv_6[4]  (.A(
        un6_next_addr_c4), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \next_addr[4]_net_1 ), .Y(\o_TPSRAM_RADDR_sv_6[4]_net_1 ));
    SLE \next_data[1]  (.D(\next_data_s[1] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[1]_net_1 ));
    GND GND (.Y(GND_net_1));
    ARI1 #( .INIT(20'h45500) )  \next_data_cry_cy[0]  (.A(VCC_net_1), 
        .B(\state_tpsram_access[0]_net_1 ), .C(GND_net_1), .D(
        GND_net_1), .FCI(VCC_net_1), .S(), .Y(), .FCO(next_data_cry_cy)
        );
    CFG4 #( .INIT(16'h7BDE) )  un1_i_TPSRAM_RD_sv_NE_2 (.A(
        \expected_data[5]_net_1 ), .B(\expected_data[4]_net_1 ), .C(
        TPSRAM_0_RD[5]), .D(TPSRAM_0_RD[4]), .Y(
        un1_i_TPSRAM_RD_sv_NE_2_net_1));
    SLE \counter[4]  (.D(\counter_s[4] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[4]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[0]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[0]_net_1 ), .Y(
        \o_TPSRAM_WD_3[0]_net_1 ));
    CFG3 #( .INIT(8'hE0) )  \state_tpsram_access_ns_a3[5]  (.A(
        o_TPSRAM_WEN8_net_1), .B(un1_i_TPSRAM_RD_sv_NE_net_1), .C(
        \state_tpsram_access[4]_net_1 ), .Y(
        \state_tpsram_access_ns_a3[5]_net_1 ));
    SLE \counter[10]  (.D(\counter_s[10] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[10]_net_1 ));
    SLE \o_TPSRAM_WADDR_sv[5]  (.D(\o_TPSRAM_WADDR_sv_3[5]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[5]));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNIVAGL5[3]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[3]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[2] ), .S(\expected_data_s[3] ), .Y(), .FCO(
        \expected_data_cry[3] ));
    SLE \counter[13]  (.D(\counter_s[13] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[13]_net_1 ));
    SLE \next_addr[1]  (.D(\next_addr_6[1]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[2]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[2]_net_1 ), .Y(
        \o_TPSRAM_WD_3[2]_net_1 ));
    SLE \counter[12]  (.D(\counter_s[12] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[12]_net_1 ));
    ARI1 #( .INIT(20'h45500) )  \counter_cry_cy[0]  (.A(VCC_net_1), .B(
        \state_tpsram_access[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), 
        .FCI(VCC_net_1), .S(), .Y(), .FCO(counter_cry_cy));
    SLE \o_TPSRAM_WD[5]  (.D(\o_TPSRAM_WD_3[5]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[5]));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNIQ13R6[4]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[4]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[3] ), .S(\expected_data_s[4] ), .Y(), .FCO(
        \expected_data_cry[4] ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[7]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[7]_net_1 ), .Y(
        \o_TPSRAM_WD_3[7]_net_1 ));
    CFG2 #( .INIT(4'h2) )  \o_TPSRAM_RADDR_sv_6[0]  (.A(
        o_TPSRAM_WEN8_RNITP5V_Y), .B(\next_addr[0]_net_1 ), .Y(
        \o_TPSRAM_RADDR_sv_6[0]_net_1 ));
    ARI1 #( .INIT(20'h4002A) )  \expected_data_RNIKCO42[0]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\expected_data[0]_net_1 ), 
        .C(o_TPSRAM_WEN8_net_1), .D(\state_tpsram_access[2]_net_1 ), 
        .FCI(expected_data_cry_cy), .S(\expected_data_s[0] ), .Y(), 
        .FCO(\expected_data_cry[0] ));
    CFG2 #( .INIT(4'h8) )  un15_0_a3 (.A(o_TPSRAM_WEN8_net_1), .B(
        \state_tpsram_access[2]_net_1 ), .Y(
        \state_tpsram_access_ns[3] ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[5]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[5]_net_1 ), .Y(
        \o_TPSRAM_WD_3[5]_net_1 ));
    SLE \counter[15]  (.D(\counter_s[15]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(countere), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\counter[15]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[3]  (.A(VCC_net_1), .B(
        \next_data[3]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[2]_net_1 ), .S(
        \next_data_s[3] ), .Y(), .FCO(\next_data_cry[3]_net_1 ));
    VCC VCC (.Y(VCC_net_1));
    CFG2 #( .INIT(4'h4) )  o_TPSRAM_WEN_RNO (.A(o_TPSRAM_WEN8_net_1), 
        .B(\state_tpsram_access[2]_net_1 ), .Y(N_90_i));
    CFG4 #( .INIT(16'h8000) )  un2_flag_1ms_11 (.A(\counter[8]_net_1 ), 
        .B(\counter[7]_net_1 ), .C(\counter[5]_net_1 ), .D(
        \counter[3]_net_1 ), .Y(un2_flag_1ms_11_net_1));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNI5LTF4[2]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[2]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[1] ), .S(\expected_data_s[2] ), .Y(), .FCO(
        \expected_data_cry[2] ));
    SLE \counter[1]  (.D(\counter_s[1] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[1]_net_1 ));
    SLE \o_TPSRAM_RADDR_sv[4]  (.D(\o_TPSRAM_RADDR_sv_6[4]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[4]));
    SLE \next_data[3]  (.D(\next_data_s[3] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[3]_net_1 ));
    SLE \expected_data[6]  (.D(\expected_data_s[6] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[6]_net_1 ));
    CFG3 #( .INIT(8'h80) )  un6_next_addr_ac0_5 (.A(
        \next_addr[2]_net_1 ), .B(o_TPSRAM_WEN8_2_net_1), .C(
        \next_addr[3]_net_1 ), .Y(un6_next_addr_c4));
    SLE o_TPSRAM_WEN (.D(N_90_i), .CLK(demo_0_FAB_CCC_GL0), .EN(
        N_103_i), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WEN));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[0]  (.A(VCC_net_1), .B(
        \counter[0]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(counter_cry_cy), .S(\counter_s[0] ), .Y(), 
        .FCO(\counter_cry[0]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[10]  (.A(VCC_net_1), .B(
        \counter[10]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[9]_net_1 ), .S(\counter_s[10] ), 
        .Y(), .FCO(\counter_cry[10]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[4]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[4]_net_1 ), .Y(
        \o_TPSRAM_WD_3[4]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  un2_flag_1ms (.A(un2_flag_1ms_11_net_1), 
        .B(un2_flag_1ms_10_net_1), .C(un2_flag_1ms_9_net_1), .D(
        un2_flag_1ms_8_net_1), .Y(N_46));
    SLE \counter[5]  (.D(\counter_s[5] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[5]_net_1 ));
    CFG4 #( .INIT(16'h48C0) )  \o_TPSRAM_RADDR_sv_6[5]  (.A(
        un6_next_addr_c4), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \next_addr[5]_net_1 ), .D(\next_addr[4]_net_1 ), .Y(
        \o_TPSRAM_RADDR_sv_6[5]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_s[7]  (.A(VCC_net_1), .B(
        \next_data[7]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[6]_net_1 ), .S(
        \next_data_s[7]_net_1 ), .Y(), .FCO());
    CFG2 #( .INIT(4'h1) )  un1_state_tpsram_access_2_0_a3 (.A(
        \state_tpsram_access[1]_net_1 ), .B(
        \state_tpsram_access[5]_net_1 ), .Y(
        un1_state_tpsram_access_2_0_a3_net_1));
    SLE \next_data[7]  (.D(\next_data_s[7]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(next_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_data[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[4]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[4]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[4]_net_1 ));
    CFG3 #( .INIT(8'h75) )  un1_i_TPSRAM_RD_sv_NE_RNI0N1L1 (.A(
        o_TPSRAM_WEN8_RNITP5V_Y), .B(un1_i_TPSRAM_RD_sv_NE_net_1), .C(
        \state_tpsram_access[4]_net_1 ), .Y(expected_datae));
    SLE \expected_data[2]  (.D(\expected_data_s[2] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[2]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[12]  (.A(VCC_net_1), .B(
        \counter[12]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[11]_net_1 ), .S(\counter_s[12] ), 
        .Y(), .FCO(\counter_cry[12]_net_1 ));
    SLE \next_data[6]  (.D(\next_data_s[6] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[6]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[2]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[2]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[0]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[0]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[0]_net_1 ));
    CFG3 #( .INIT(8'h60) )  \o_TPSRAM_RADDR_sv_6[1]  (.A(
        \next_addr[1]_net_1 ), .B(\next_addr[0]_net_1 ), .C(
        o_TPSRAM_WEN8_RNITP5V_Y), .Y(\o_TPSRAM_RADDR_sv_6[1]_net_1 ));
    ARI1 #( .INIT(20'h41500) )  o_TPSRAM_WEN8_RNITP5V (.A(VCC_net_1), 
        .B(\state_tpsram_access[0]_net_1 ), .C(
        \state_tpsram_access[2]_net_1 ), .D(o_TPSRAM_WEN8_net_1), .FCI(
        VCC_net_1), .S(), .Y(o_TPSRAM_WEN8_RNITP5V_Y), .FCO(
        expected_data_cry_cy));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[1]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[1]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[1]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[5]  (.A(VCC_net_1), .B(
        \next_data[5]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[4]_net_1 ), .S(
        \next_data_s[5] ), .Y(), .FCO(\next_data_cry[5]_net_1 ));
    SLE \state_tpsram_access[4]  (.D(\state_tpsram_access_ns[4]_net_1 )
        , .CLK(demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[4]_net_1 ));
    CFG4 #( .INIT(16'h48C0) )  \o_TPSRAM_RADDR_sv_6[3]  (.A(
        o_TPSRAM_WEN8_2_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \next_addr[3]_net_1 ), .D(\next_addr[2]_net_1 ), .Y(
        \o_TPSRAM_RADDR_sv_6[3]_net_1 ));
    SLE \o_TPSRAM_WADDR_sv[4]  (.D(\o_TPSRAM_WADDR_sv_3[4]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[4]));
    CFG3 #( .INIT(8'h06) )  \next_addr_6[2]  (.A(\next_addr[2]_net_1 ), 
        .B(o_TPSRAM_WEN8_2_net_1), .C(un1_state_tpsram_access_10), .Y(
        \next_addr_6[2]_net_1 ));
    CFG4 #( .INIT(16'h7BDE) )  un1_i_TPSRAM_RD_sv_NE_1 (.A(
        \expected_data[3]_net_1 ), .B(\expected_data[2]_net_1 ), .C(
        TPSRAM_0_RD[3]), .D(TPSRAM_0_RD[2]), .Y(
        un1_i_TPSRAM_RD_sv_NE_1_net_1));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[14]  (.A(VCC_net_1), .B(
        \counter[14]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[13]_net_1 ), .S(\counter_s[14] ), 
        .Y(), .FCO(\counter_cry[14]_net_1 ));
    SLE o_reset_n (.D(\state_tpsram_access[0]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_7_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(Ram_intferface_0_o_reset_n)
        );
    SLE \counter[14]  (.D(\counter_s[14] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[14]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[1]  (.A(VCC_net_1), .B(
        \counter[1]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[0]_net_1 ), .S(\counter_s[1] ), 
        .Y(), .FCO(\counter_cry[1]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[11]  (.A(VCC_net_1), .B(
        \counter[11]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[10]_net_1 ), .S(\counter_s[11] ), 
        .Y(), .FCO(\counter_cry[11]_net_1 ));
    CFG4 #( .INIT(16'hA3A0) )  \state_tpsram_access_RNO[2]  (.A(N_46), 
        .B(o_TPSRAM_WEN8_net_1), .C(\state_tpsram_access[1]_net_1 ), 
        .D(\state_tpsram_access[2]_net_1 ), .Y(N_76_i));
    SLE \next_data[0]  (.D(\next_data_s[0] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[0]_net_1 ));
    CFG2 #( .INIT(4'h1) )  \next_addr_6[0]  (.A(
        un1_state_tpsram_access_10), .B(\next_addr[0]_net_1 ), .Y(
        \next_addr_6[0]_net_1 ));
    CFG3 #( .INIT(8'h8F) )  un1_state_tpsram_access_10_0 (.A(
        \state_tpsram_access[4]_net_1 ), .B(o_TPSRAM_WEN8_net_1), .C(
        o_TPSRAM_WEN8_RNITP5V_Y), .Y(un1_state_tpsram_access_10));
    CFG2 #( .INIT(4'h8) )  o_TPSRAM_WEN8_2 (.A(\next_addr[0]_net_1 ), 
        .B(\next_addr[1]_net_1 ), .Y(o_TPSRAM_WEN8_2_net_1));
    SLE \state_tpsram_access[0]  (.D(GND_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(GND_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[0]_net_1 ));
    SLE \next_addr[2]  (.D(\next_addr_6[2]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[2]_net_1 ));
    SLE \expected_data[3]  (.D(\expected_data_s[3] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[3]_net_1 ));
    SLE \state_tpsram_access[5]  (.D(VCC_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(\state_tpsram_access_ns_a3[5]_net_1 ), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[5]_net_1 ));
    CFG4 #( .INIT(16'h060C) )  \next_addr_6[3]  (.A(
        \next_addr[2]_net_1 ), .B(\next_addr[3]_net_1 ), .C(
        un1_state_tpsram_access_10), .D(o_TPSRAM_WEN8_2_net_1), .Y(
        \next_addr_6[3]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  un2_flag_1ms_10 (.A(\counter[14]_net_1 )
        , .B(\counter[13]_net_1 ), .C(\counter[1]_net_1 ), .D(
        \counter[0]_net_1 ), .Y(un2_flag_1ms_10_net_1));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[6]  (.A(VCC_net_1), .B(
        \counter[6]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[5]_net_1 ), .S(\counter_s[6] ), 
        .Y(), .FCO(\counter_cry[6]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_s[15]  (.A(VCC_net_1), .B(
        \counter[15]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[14]_net_1 ), .S(
        \counter_s[15]_net_1 ), .Y(), .FCO());
    CFG3 #( .INIT(8'hDC) )  \un1_state_tpsram_access_4_0[0]  (.A(
        o_TPSRAM_WEN8_net_1), .B(\state_tpsram_access_ns[3] ), .C(
        \state_tpsram_access[4]_net_1 ), .Y(
        \un1_state_tpsram_access_4[0] ));
    SLE \state_tpsram_access[1]  (.D(\state_tpsram_access_ns[1]_net_1 )
        , .CLK(demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[1]_net_1 ));
    SLE \o_TPSRAM_WD[3]  (.D(\o_TPSRAM_WD_3[3]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[3]));
    CFG2 #( .INIT(4'hE) )  \state_tpsram_access_RNIGRPG[2]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(
        \state_tpsram_access[2]_net_1 ), .Y(N_103_i));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[5]  (.A(VCC_net_1), .B(
        \counter[5]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[4]_net_1 ), .S(\counter_s[5] ), 
        .Y(), .FCO(\counter_cry[5]_net_1 ));
    SLE \o_TPSRAM_WD[1]  (.D(\o_TPSRAM_WD_3[1]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[1]));
    CFG3 #( .INIT(8'h12) )  \next_addr_6[1]  (.A(\next_addr[0]_net_1 ), 
        .B(un1_state_tpsram_access_10), .C(\next_addr[1]_net_1 ), .Y(
        \next_addr_6[1]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[4]  (.A(VCC_net_1), .B(
        \next_data[4]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[3]_net_1 ), .S(
        \next_data_s[4] ), .Y(), .FCO(\next_data_cry[4]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[8]  (.A(VCC_net_1), .B(
        \counter[8]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[7]_net_1 ), .S(\counter_s[8] ), 
        .Y(), .FCO(\counter_cry[8]_net_1 ));
    SLE \counter[7]  (.D(\counter_s[7] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[7]_net_1 ));
    SLE \next_addr[5]  (.D(\next_addr_6[5]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[5]_net_1 ));
    CFG3 #( .INIT(8'hFE) )  un15_0 (.A(\state_tpsram_access[0]_net_1 ), 
        .B(\state_tpsram_access_ns[3] ), .C(
        \state_tpsram_access[4]_net_1 ), .Y(un15_0_net_1));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WD_3[6]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_data[6]_net_1 ), .Y(
        \o_TPSRAM_WD_3[6]_net_1 ));
    SLE \next_data[2]  (.D(\next_data_s[2] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(next_datae), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1)
        , .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \next_data[2]_net_1 ));
    CFG4 #( .INIT(16'h7BDE) )  un1_i_TPSRAM_RD_sv_NE_3 (.A(
        \expected_data[7]_net_1 ), .B(\expected_data[6]_net_1 ), .C(
        TPSRAM_0_RD[7]), .D(TPSRAM_0_RD[6]), .Y(
        un1_i_TPSRAM_RD_sv_NE_3_net_1));
    SLE \o_TPSRAM_RADDR_sv[0]  (.D(\o_TPSRAM_RADDR_sv_6[0]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[0]));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[7]  (.A(VCC_net_1), .B(
        \counter[7]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[6]_net_1 ), .S(\counter_s[7] ), 
        .Y(), .FCO(\counter_cry[7]_net_1 ));
    CFG4 #( .INIT(16'h7BDE) )  un1_i_TPSRAM_RD_sv_NE_0 (.A(
        \expected_data[1]_net_1 ), .B(\expected_data[0]_net_1 ), .C(
        TPSRAM_0_RD[1]), .D(TPSRAM_0_RD[0]), .Y(
        un1_i_TPSRAM_RD_sv_NE_0_net_1));
    SLE o_TPSRAM_REN (.D(\un1_state_tpsram_access_4[0] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un15_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_REN));
    SLE \expected_data[7]  (.D(\expected_data_s[7] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[7]_net_1 ));
    CFG4 #( .INIT(16'hFFFE) )  un1_i_TPSRAM_RD_sv_NE (.A(
        un1_i_TPSRAM_RD_sv_NE_3_net_1), .B(
        un1_i_TPSRAM_RD_sv_NE_2_net_1), .C(
        un1_i_TPSRAM_RD_sv_NE_1_net_1), .D(
        un1_i_TPSRAM_RD_sv_NE_0_net_1), .Y(un1_i_TPSRAM_RD_sv_NE_net_1)
        );
    ARI1 #( .INIT(20'h42200) )  \counter_cry[9]  (.A(VCC_net_1), .B(
        \counter[9]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[8]_net_1 ), .S(\counter_s[9] ), 
        .Y(), .FCO(\counter_cry[9]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[1]  (.A(VCC_net_1), .B(
        \next_data[1]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[0]_net_1 ), .S(
        \next_data_s[1] ), .Y(), .FCO(\next_data_cry[1]_net_1 ));
    CFG4 #( .INIT(16'h006A) )  \next_addr_6[5]  (.A(
        \next_addr[5]_net_1 ), .B(\next_addr[4]_net_1 ), .C(
        un6_next_addr_c4), .D(un1_state_tpsram_access_10), .Y(
        \next_addr_6[5]_net_1 ));
    CFG3 #( .INIT(8'h48) )  \o_TPSRAM_RADDR_sv_6[2]  (.A(
        o_TPSRAM_WEN8_2_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \next_addr[2]_net_1 ), .Y(\o_TPSRAM_RADDR_sv_6[2]_net_1 ));
    SLE \o_TPSRAM_WD[2]  (.D(\o_TPSRAM_WD_3[2]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WD[2]));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNIJI869[6]  (.A(
        VCC_net_1), .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(
        \expected_data[6]_net_1 ), .D(GND_net_1), .FCI(
        \expected_data_cry[5] ), .S(\expected_data_s[6] ), .Y(), .FCO(
        \expected_data_cry[6] ));
    SLE \expected_data[5]  (.D(\expected_data_s[5] ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(expected_datae), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(\expected_data[5]_net_1 ));
    SLE \o_TPSRAM_RADDR_sv[1]  (.D(\o_TPSRAM_RADDR_sv_6[1]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[1]));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[2]  (.A(VCC_net_1), .B(
        \counter[2]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[1]_net_1 ), .S(\counter_s[2] ), 
        .Y(), .FCO(\counter_cry[2]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[2]  (.A(VCC_net_1), .B(
        \next_data[2]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(\next_data_cry[1]_net_1 ), .S(
        \next_data_s[2] ), .Y(), .FCO(\next_data_cry[2]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[5]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[5]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[5]_net_1 ));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[4]  (.A(VCC_net_1), .B(
        \counter[4]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[3]_net_1 ), .S(\counter_s[4] ), 
        .Y(), .FCO(\counter_cry[4]_net_1 ));
    SLE \counter[9]  (.D(\counter_s[9] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[9]_net_1 ));
    ARI1 #( .INIT(20'h48800) )  \expected_data_RNO[7]  (.A(VCC_net_1), 
        .B(o_TPSRAM_WEN8_RNITP5V_Y), .C(\expected_data[7]_net_1 ), .D(
        GND_net_1), .FCI(\expected_data_cry[6] ), .S(
        \expected_data_s[7] ), .Y(), .FCO());
    SLE \state_tpsram_access[3]  (.D(\state_tpsram_access_ns[3] ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \state_tpsram_access[3]_net_1 ));
    SLE \o_TPSRAM_RADDR_sv[2]  (.D(\o_TPSRAM_RADDR_sv_6[2]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[2]));
    CFG2 #( .INIT(4'hE) )  \state_tpsram_access_RNIHSPG[1]  (.A(
        \state_tpsram_access[2]_net_1 ), .B(
        \state_tpsram_access[1]_net_1 ), .Y(countere));
    SLE \o_TPSRAM_RADDR_sv[3]  (.D(\o_TPSRAM_RADDR_sv_6[3]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(
        un1_state_tpsram_access_9_0_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_RADDR_sv[3]));
    ARI1 #( .INIT(20'h42200) )  \counter_cry[13]  (.A(VCC_net_1), .B(
        \counter[13]_net_1 ), .C(\state_tpsram_access[2]_net_1 ), .D(
        GND_net_1), .FCI(\counter_cry[12]_net_1 ), .S(\counter_s[13] ), 
        .Y(), .FCO(\counter_cry[13]_net_1 ));
    SLE \counter[8]  (.D(\counter_s[8] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[8]_net_1 ));
    SLE \o_TPSRAM_WADDR_sv[0]  (.D(\o_TPSRAM_WADDR_sv_3[0]_net_1 ), 
        .CLK(demo_0_FAB_CCC_GL0), .EN(N_103_i), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        Ram_intferface_0_o_TPSRAM_WADDR_sv[0]));
    ARI1 #( .INIT(20'h42200) )  \next_data_cry[0]  (.A(VCC_net_1), .B(
        \next_data[0]_net_1 ), .C(\state_tpsram_access[0]_net_1 ), .D(
        GND_net_1), .FCI(next_data_cry_cy), .S(\next_data_s[0] ), .Y(), 
        .FCO(\next_data_cry[0]_net_1 ));
    CFG2 #( .INIT(4'h1) )  o_TPSRAM_WEN8_1 (.A(\next_addr[4]_net_1 ), 
        .B(\next_addr[3]_net_1 ), .Y(o_TPSRAM_WEN8_1_net_1));
    CFG3 #( .INIT(8'hCE) )  o_TPSRAM_WEN8_RNITP5V_0 (.A(
        \state_tpsram_access[2]_net_1 ), .B(
        \state_tpsram_access[0]_net_1 ), .C(o_TPSRAM_WEN8_net_1), .Y(
        next_datae));
    CFG2 #( .INIT(4'h4) )  \o_TPSRAM_WADDR_sv_3[3]  (.A(
        \state_tpsram_access[0]_net_1 ), .B(\next_addr[3]_net_1 ), .Y(
        \o_TPSRAM_WADDR_sv_3[3]_net_1 ));
    CFG3 #( .INIT(8'h14) )  \next_addr_6[4]  (.A(
        un1_state_tpsram_access_10), .B(\next_addr[4]_net_1 ), .C(
        un6_next_addr_c4), .Y(\next_addr_6[4]_net_1 ));
    SLE \counter[0]  (.D(\counter_s[0] ), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(countere), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        \counter[0]_net_1 ));
    SLE \next_addr[3]  (.D(\next_addr_6[3]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(un1_state_tpsram_access_2_0_a3_net_1), 
        .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1)
        , .SD(GND_net_1), .LAT(GND_net_1), .Q(\next_addr[3]_net_1 ));
    
endmodule


module Dev_Restart_after_ISP_blk_TPSRAM_0_TPSRAM(
       Ram_intferface_0_o_TPSRAM_WADDR_sv,
       Ram_intferface_0_o_TPSRAM_WD,
       Ram_intferface_0_o_TPSRAM_RADDR_sv,
       TPSRAM_0_RD,
       Ram_intferface_0_o_TPSRAM_WEN,
       Ram_intferface_0_o_TPSRAM_REN,
       demo_0_FAB_CCC_GL0
    );
input  [5:0] Ram_intferface_0_o_TPSRAM_WADDR_sv;
input  [7:0] Ram_intferface_0_o_TPSRAM_WD;
input  [5:0] Ram_intferface_0_o_TPSRAM_RADDR_sv;
output [7:0] TPSRAM_0_RD;
input  Ram_intferface_0_o_TPSRAM_WEN;
input  Ram_intferface_0_o_TPSRAM_REN;
input  demo_0_FAB_CCC_GL0;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    RAM1K18 Dev_Restart_after_ISP_blk_TPSRAM_0_TPSRAM_R0C0 (.A_DOUT({
        nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7, nc8, nc9, 
        TPSRAM_0_RD[7], TPSRAM_0_RD[6], TPSRAM_0_RD[5], TPSRAM_0_RD[4], 
        TPSRAM_0_RD[3], TPSRAM_0_RD[2], TPSRAM_0_RD[1], TPSRAM_0_RD[0]})
        , .B_DOUT({nc10, nc11, nc12, nc13, nc14, nc15, nc16, nc17, 
        nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, nc26, nc27}), 
        .BUSY(), .A_CLK(demo_0_FAB_CCC_GL0), .A_DOUT_CLK(VCC_net_1), 
        .A_ARST_N(VCC_net_1), .A_DOUT_EN(VCC_net_1), .A_BLK({
        Ram_intferface_0_o_TPSRAM_REN, VCC_net_1, VCC_net_1}), 
        .A_DOUT_ARST_N(VCC_net_1), .A_DOUT_SRST_N(VCC_net_1), .A_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .A_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[5], 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[4], 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[3], 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[2], 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[1], 
        Ram_intferface_0_o_TPSRAM_RADDR_sv[0], GND_net_1, GND_net_1, 
        GND_net_1}), .A_WEN({GND_net_1, GND_net_1}), .B_CLK(
        demo_0_FAB_CCC_GL0), .B_DOUT_CLK(VCC_net_1), .B_ARST_N(
        VCC_net_1), .B_DOUT_EN(VCC_net_1), .B_BLK({
        Ram_intferface_0_o_TPSRAM_WEN, VCC_net_1, VCC_net_1}), 
        .B_DOUT_ARST_N(GND_net_1), .B_DOUT_SRST_N(VCC_net_1), .B_DIN({
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Ram_intferface_0_o_TPSRAM_WD[7], 
        Ram_intferface_0_o_TPSRAM_WD[6], 
        Ram_intferface_0_o_TPSRAM_WD[5], 
        Ram_intferface_0_o_TPSRAM_WD[4], 
        Ram_intferface_0_o_TPSRAM_WD[3], 
        Ram_intferface_0_o_TPSRAM_WD[2], 
        Ram_intferface_0_o_TPSRAM_WD[1], 
        Ram_intferface_0_o_TPSRAM_WD[0]}), .B_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[5], 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[4], 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[3], 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[2], 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[1], 
        Ram_intferface_0_o_TPSRAM_WADDR_sv[0], GND_net_1, GND_net_1, 
        GND_net_1}), .B_WEN({GND_net_1, VCC_net_1}), .A_EN(VCC_net_1), 
        .A_DOUT_LAT(VCC_net_1), .A_WIDTH({GND_net_1, VCC_net_1, 
        VCC_net_1}), .A_WMODE(GND_net_1), .B_EN(VCC_net_1), 
        .B_DOUT_LAT(VCC_net_1), .B_WIDTH({GND_net_1, VCC_net_1, 
        VCC_net_1}), .B_WMODE(GND_net_1), .SII_LOCK(GND_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module Dev_Restart_after_ISP_blk_TAMPER2_0_TAMPER2(
       Ram_intferface_0_o_reset_n
    );
input  Ram_intferface_0_o_reset_n;

    wire VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    TAMPER TAMPER_INST (.JTAG_ACTIVE(), .LOCK_TAMPER_DETECT(), 
        .MESH_SHORT_ERROR(), .CLK_ERROR(), .DETECT_CATEGORY({nc0, nc1, 
        nc2, nc3}), .DETECT_ATTEMPT(), .DETECT_FAIL(), .DIGEST_ERROR(), 
        .POWERUP_DIGEST_ERROR(), .SC_ROM_DIGEST_ERROR(), 
        .TAMPER_CHANGE_STROBE(), .LOCKDOWN_ALL_N(VCC_net_1), 
        .DISABLE_ALL_IOS_N(VCC_net_1), .RESET_N(
        Ram_intferface_0_o_reset_n), .ZEROIZE_N(VCC_net_1));
    
endmodule


module Dev_Restart_after_ISP_blk(
       demo_0_POWER_ON_RESET_N,
       demo_0_FAB_CCC_GL0
    );
input  demo_0_POWER_ON_RESET_N;
input  demo_0_FAB_CCC_GL0;

    wire \TPSRAM_0_RD[0] , \TPSRAM_0_RD[1] , \TPSRAM_0_RD[2] , 
        \TPSRAM_0_RD[3] , \TPSRAM_0_RD[4] , \TPSRAM_0_RD[5] , 
        \TPSRAM_0_RD[6] , \TPSRAM_0_RD[7] , 
        \Ram_intferface_0_o_TPSRAM_WD[0] , 
        \Ram_intferface_0_o_TPSRAM_WD[1] , 
        \Ram_intferface_0_o_TPSRAM_WD[2] , 
        \Ram_intferface_0_o_TPSRAM_WD[3] , 
        \Ram_intferface_0_o_TPSRAM_WD[4] , 
        \Ram_intferface_0_o_TPSRAM_WD[5] , 
        \Ram_intferface_0_o_TPSRAM_WD[6] , 
        \Ram_intferface_0_o_TPSRAM_WD[7] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[0] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[5] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[0] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[5] , 
        Ram_intferface_0_o_TPSRAM_REN, Ram_intferface_0_o_TPSRAM_WEN, 
        Ram_intferface_0_o_reset_n, GND_net_1, VCC_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    Ram_intferface Ram_intferface_0 (.TPSRAM_0_RD({\TPSRAM_0_RD[7] , 
        \TPSRAM_0_RD[6] , \TPSRAM_0_RD[5] , \TPSRAM_0_RD[4] , 
        \TPSRAM_0_RD[3] , \TPSRAM_0_RD[2] , \TPSRAM_0_RD[1] , 
        \TPSRAM_0_RD[0] }), .Ram_intferface_0_o_TPSRAM_WD({
        \Ram_intferface_0_o_TPSRAM_WD[7] , 
        \Ram_intferface_0_o_TPSRAM_WD[6] , 
        \Ram_intferface_0_o_TPSRAM_WD[5] , 
        \Ram_intferface_0_o_TPSRAM_WD[4] , 
        \Ram_intferface_0_o_TPSRAM_WD[3] , 
        \Ram_intferface_0_o_TPSRAM_WD[2] , 
        \Ram_intferface_0_o_TPSRAM_WD[1] , 
        \Ram_intferface_0_o_TPSRAM_WD[0] }), 
        .Ram_intferface_0_o_TPSRAM_RADDR_sv({
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[5] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[0] }), 
        .Ram_intferface_0_o_TPSRAM_WADDR_sv({
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[5] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[0] }), 
        .Ram_intferface_0_o_TPSRAM_REN(Ram_intferface_0_o_TPSRAM_REN), 
        .Ram_intferface_0_o_TPSRAM_WEN(Ram_intferface_0_o_TPSRAM_WEN), 
        .Ram_intferface_0_o_reset_n(Ram_intferface_0_o_reset_n), 
        .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0), 
        .demo_0_POWER_ON_RESET_N(demo_0_POWER_ON_RESET_N));
    Dev_Restart_after_ISP_blk_TPSRAM_0_TPSRAM TPSRAM_0 (
        .Ram_intferface_0_o_TPSRAM_WADDR_sv({
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[5] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_WADDR_sv[0] }), 
        .Ram_intferface_0_o_TPSRAM_WD({
        \Ram_intferface_0_o_TPSRAM_WD[7] , 
        \Ram_intferface_0_o_TPSRAM_WD[6] , 
        \Ram_intferface_0_o_TPSRAM_WD[5] , 
        \Ram_intferface_0_o_TPSRAM_WD[4] , 
        \Ram_intferface_0_o_TPSRAM_WD[3] , 
        \Ram_intferface_0_o_TPSRAM_WD[2] , 
        \Ram_intferface_0_o_TPSRAM_WD[1] , 
        \Ram_intferface_0_o_TPSRAM_WD[0] }), 
        .Ram_intferface_0_o_TPSRAM_RADDR_sv({
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[5] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[4] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[3] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[2] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[1] , 
        \Ram_intferface_0_o_TPSRAM_RADDR_sv[0] }), .TPSRAM_0_RD({
        \TPSRAM_0_RD[7] , \TPSRAM_0_RD[6] , \TPSRAM_0_RD[5] , 
        \TPSRAM_0_RD[4] , \TPSRAM_0_RD[3] , \TPSRAM_0_RD[2] , 
        \TPSRAM_0_RD[1] , \TPSRAM_0_RD[0] }), 
        .Ram_intferface_0_o_TPSRAM_WEN(Ram_intferface_0_o_TPSRAM_WEN), 
        .Ram_intferface_0_o_TPSRAM_REN(Ram_intferface_0_o_TPSRAM_REN), 
        .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0));
    Dev_Restart_after_ISP_blk_TAMPER2_0_TAMPER2 TAMPER2_0 (
        .Ram_intferface_0_o_reset_n(Ram_intferface_0_o_reset_n));
    
endmodule


module BLINK_LED(
       LED1_c,
       demo_0_FAB_CCC_GL0,
       demo_0_MSS_READY
    );
output LED1_c;
input  demo_0_FAB_CCC_GL0;
input  demo_0_MSS_READY;

    wire \counter[29]_net_1 , VCC_net_1, un2_counter_1_cry_29_S, 
        GND_net_1, \counter[30]_net_1 , un2_counter_1_cry_30_S, 
        \counter[31]_net_1 , un2_counter_1_s_31_S, \counter[14]_net_1 , 
        \counter_4[14]_net_1 , \counter[15]_net_1 , 
        un2_counter_1_cry_15_S, \counter[16]_net_1 , 
        un2_counter_1_cry_16_S, \counter[17]_net_1 , 
        \counter_4[17]_net_1 , \counter[18]_net_1 , 
        un2_counter_1_cry_18_S, \counter[19]_net_1 , 
        un2_counter_1_cry_19_S, \counter[20]_net_1 , 
        un2_counter_1_cry_20_S, \counter[21]_net_1 , 
        \counter_4[21]_net_1 , \counter[22]_net_1 , 
        \counter_4[22]_net_1 , \counter[23]_net_1 , 
        un2_counter_1_cry_23_S, \counter[24]_net_1 , 
        un2_counter_1_cry_24_S, \counter[25]_net_1 , 
        \counter_4[25]_net_1 , \counter[26]_net_1 , 
        un2_counter_1_cry_26_S, \counter[27]_net_1 , 
        un2_counter_1_cry_27_S, \counter[28]_net_1 , 
        un2_counter_1_cry_28_S, \counter[0]_net_1 , 
        \counter_4[0]_net_1 , \counter[1]_net_1 , 
        un2_counter_1_cry_1_S, \counter[2]_net_1 , 
        un2_counter_1_cry_2_S, \counter[3]_net_1 , 
        un2_counter_1_cry_3_S, \counter[4]_net_1 , 
        un2_counter_1_cry_4_S, \counter[5]_net_1 , 
        un2_counter_1_cry_5_S, \counter[6]_net_1 , 
        un2_counter_1_cry_6_S, \counter[7]_net_1 , 
        un2_counter_1_cry_7_S, \counter[8]_net_1 , 
        un2_counter_1_cry_8_S, \counter[9]_net_1 , 
        \counter_4[9]_net_1 , \counter[10]_net_1 , 
        un2_counter_1_cry_10_S, \counter[11]_net_1 , 
        \counter_4[11]_net_1 , \counter[12]_net_1 , 
        \counter_4[12]_net_1 , \counter[13]_net_1 , 
        un2_counter_1_cry_13_S, LED1_0_net_1, un2_counter_1_s_1_90_FCO, 
        un2_counter_1_cry_1_net_1, un2_counter_1_cry_2_net_1, 
        un2_counter_1_cry_3_net_1, un2_counter_1_cry_4_net_1, 
        un2_counter_1_cry_5_net_1, un2_counter_1_cry_6_net_1, 
        un2_counter_1_cry_7_net_1, un2_counter_1_cry_8_net_1, 
        un2_counter_1_cry_9_net_1, un2_counter_1_cry_9_S, 
        un2_counter_1_cry_10_net_1, un2_counter_1_cry_11_net_1, 
        un2_counter_1_cry_11_S, un2_counter_1_cry_12_net_1, 
        un2_counter_1_cry_12_S, un2_counter_1_cry_13_net_1, 
        un2_counter_1_cry_14_net_1, un2_counter_1_cry_14_S, 
        un2_counter_1_cry_15_net_1, un2_counter_1_cry_16_net_1, 
        un2_counter_1_cry_17_net_1, un2_counter_1_cry_17_S, 
        un2_counter_1_cry_18_net_1, un2_counter_1_cry_19_net_1, 
        un2_counter_1_cry_20_net_1, un2_counter_1_cry_21_net_1, 
        un2_counter_1_cry_21_S, un2_counter_1_cry_22_net_1, 
        un2_counter_1_cry_22_S, un2_counter_1_cry_23_net_1, 
        un2_counter_1_cry_24_net_1, un2_counter_1_cry_25_net_1, 
        un2_counter_1_cry_25_S, un2_counter_1_cry_26_net_1, 
        un2_counter_1_cry_27_net_1, un2_counter_1_cry_28_net_1, 
        un2_counter_1_cry_29_net_1, un2_counter_1_cry_30_net_1, 
        counter12_18_net_1, counter12_17_net_1, counter12_16_net_1, 
        counter12_15_net_1, counter12_14_net_1, counter12_13_net_1, 
        counter11_19_net_1, counter11_18_net_1, counter11_17_net_1, 
        counter11_16_net_1, counter11_15_net_1, counter11_14_net_1, 
        counter11_13_net_1, counter11_20_net_1, counter12_19_net_1, 
        counter12_24_net_1, counter11_25_net_1, counter11_24_net_1, 
        counter12_net_1;
    
    CFG2 #( .INIT(4'h4) )  \counter_4[25]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_25_S), .Y(\counter_4[25]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_20 (.A(VCC_net_1), 
        .B(\counter[20]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_19_net_1), .S(un2_counter_1_cry_20_S), .Y(), 
        .FCO(un2_counter_1_cry_20_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_13 (.A(VCC_net_1), 
        .B(\counter[13]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_12_net_1), .S(un2_counter_1_cry_13_S), .Y(), 
        .FCO(un2_counter_1_cry_13_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_1 (.A(VCC_net_1), .B(
        \counter[1]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_s_1_90_FCO), .S(un2_counter_1_cry_1_S), .Y(), 
        .FCO(un2_counter_1_cry_1_net_1));
    SLE \counter[24]  (.D(un2_counter_1_cry_24_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[24]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_4 (.A(VCC_net_1), .B(
        \counter[4]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_3_net_1), .S(un2_counter_1_cry_4_S), .Y(), 
        .FCO(un2_counter_1_cry_4_net_1));
    SLE \counter[17]  (.D(\counter_4[17]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[17]_net_1 ));
    CFG4 #( .INIT(16'h4000) )  counter12_19 (.A(\counter[23]_net_1 ), 
        .B(\counter[11]_net_1 ), .C(\counter[9]_net_1 ), .D(
        counter12_13_net_1), .Y(counter12_19_net_1));
    SLE \counter[2]  (.D(un2_counter_1_cry_2_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[2]_net_1 ));
    SLE \counter[7]  (.D(un2_counter_1_cry_7_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[7]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \counter_4[22]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_22_S), .Y(\counter_4[22]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \counter_4[11]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_11_S), .Y(\counter_4[11]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_28 (.A(VCC_net_1), 
        .B(\counter[28]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_27_net_1), .S(un2_counter_1_cry_28_S), .Y(), 
        .FCO(un2_counter_1_cry_28_net_1));
    CFG2 #( .INIT(4'h4) )  \counter_4[9]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_9_S), .Y(\counter_4[9]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter12_15 (.A(\counter[24]_net_1 ), 
        .B(\counter[20]_net_1 ), .C(\counter[16]_net_1 ), .D(
        \counter[13]_net_1 ), .Y(counter12_15_net_1));
    SLE \counter[6]  (.D(un2_counter_1_cry_6_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[6]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_s_31 (.A(VCC_net_1), .B(
        \counter[31]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_30_net_1), .S(un2_counter_1_s_31_S), .Y(), 
        .FCO());
    SLE LED1 (.D(LED1_0_net_1), .CLK(demo_0_FAB_CCC_GL0), .EN(
        VCC_net_1), .ALn(demo_0_MSS_READY), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(LED1_c));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_15 (.A(VCC_net_1), 
        .B(\counter[15]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_14_net_1), .S(un2_counter_1_cry_15_S), .Y(), 
        .FCO(un2_counter_1_cry_15_net_1));
    CFG4 #( .INIT(16'h0001) )  counter11_17 (.A(\counter[5]_net_1 ), 
        .B(\counter[4]_net_1 ), .C(\counter[3]_net_1 ), .D(
        \counter[2]_net_1 ), .Y(counter11_17_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE \counter[8]  (.D(un2_counter_1_cry_8_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[8]_net_1 ));
    SLE \counter[22]  (.D(\counter_4[22]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[22]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter11_16 (.A(\counter[25]_net_1 ), 
        .B(\counter[22]_net_1 ), .C(\counter[1]_net_1 ), .D(
        \counter[0]_net_1 ), .Y(counter11_16_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_14 (.A(VCC_net_1), 
        .B(\counter[14]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_13_net_1), .S(un2_counter_1_cry_14_S), .Y(), 
        .FCO(un2_counter_1_cry_14_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_5 (.A(VCC_net_1), .B(
        \counter[5]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_4_net_1), .S(un2_counter_1_cry_5_S), .Y(), 
        .FCO(un2_counter_1_cry_5_net_1));
    SLE \counter[16]  (.D(un2_counter_1_cry_16_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[16]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_s_1_90 (.A(VCC_net_1), 
        .B(\counter[0]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        VCC_net_1), .S(), .Y(), .FCO(un2_counter_1_s_1_90_FCO));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_8 (.A(VCC_net_1), .B(
        \counter[8]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_7_net_1), .S(un2_counter_1_cry_8_S), .Y(), 
        .FCO(un2_counter_1_cry_8_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_19 (.A(VCC_net_1), 
        .B(\counter[19]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_18_net_1), .S(un2_counter_1_cry_19_S), .Y(), 
        .FCO(un2_counter_1_cry_19_net_1));
    SLE \counter[15]  (.D(un2_counter_1_cry_15_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[15]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_9 (.A(VCC_net_1), .B(
        \counter[9]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_8_net_1), .S(un2_counter_1_cry_9_S), .Y(), 
        .FCO(un2_counter_1_cry_9_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_27 (.A(VCC_net_1), 
        .B(\counter[27]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_26_net_1), .S(un2_counter_1_cry_27_S), .Y(), 
        .FCO(un2_counter_1_cry_27_net_1));
    SLE \counter[29]  (.D(un2_counter_1_cry_29_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[29]_net_1 ));
    CFG4 #( .INIT(16'h0008) )  counter12_14 (.A(\counter[25]_net_1 ), 
        .B(\counter[22]_net_1 ), .C(\counter[10]_net_1 ), .D(
        \counter[8]_net_1 ), .Y(counter12_14_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_21 (.A(VCC_net_1), 
        .B(\counter[21]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_20_net_1), .S(un2_counter_1_cry_21_S), .Y(), 
        .FCO(un2_counter_1_cry_21_net_1));
    CFG4 #( .INIT(16'h8000) )  counter11_13 (.A(\counter[13]_net_1 ), 
        .B(\counter[11]_net_1 ), .C(\counter[10]_net_1 ), .D(
        \counter[8]_net_1 ), .Y(counter11_13_net_1));
    SLE \counter[14]  (.D(\counter_4[14]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[14]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_22 (.A(VCC_net_1), 
        .B(\counter[22]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_21_net_1), .S(un2_counter_1_cry_22_S), .Y(), 
        .FCO(un2_counter_1_cry_22_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_10 (.A(VCC_net_1), 
        .B(\counter[10]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_9_net_1), .S(un2_counter_1_cry_10_S), .Y(), 
        .FCO(un2_counter_1_cry_10_net_1));
    CFG3 #( .INIT(8'h6A) )  LED1_0 (.A(LED1_c), .B(counter11_25_net_1), 
        .C(counter11_24_net_1), .Y(LED1_0_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_26 (.A(VCC_net_1), 
        .B(\counter[26]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_25_net_1), .S(un2_counter_1_cry_26_S), .Y(), 
        .FCO(un2_counter_1_cry_26_net_1));
    SLE \counter[21]  (.D(\counter_4[21]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[21]_net_1 ));
    GND GND (.Y(GND_net_1));
    SLE \counter[4]  (.D(un2_counter_1_cry_4_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[4]_net_1 ));
    SLE \counter[28]  (.D(un2_counter_1_cry_28_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[28]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter11_18 (.A(\counter[18]_net_1 ), 
        .B(\counter[15]_net_1 ), .C(\counter[7]_net_1 ), .D(
        \counter[6]_net_1 ), .Y(counter11_18_net_1));
    SLE \counter[5]  (.D(un2_counter_1_cry_5_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[5]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_3 (.A(VCC_net_1), .B(
        \counter[3]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_2_net_1), .S(un2_counter_1_cry_3_S), .Y(), 
        .FCO(un2_counter_1_cry_3_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_18 (.A(VCC_net_1), 
        .B(\counter[18]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_17_net_1), .S(un2_counter_1_cry_18_S), .Y(), 
        .FCO(un2_counter_1_cry_18_net_1));
    SLE \counter[31]  (.D(un2_counter_1_s_31_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[31]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  counter12 (.A(counter12_14_net_1), .B(
        counter12_15_net_1), .C(counter12_24_net_1), .D(
        counter12_19_net_1), .Y(counter12_net_1));
    CFG4 #( .INIT(16'h8000) )  counter11_25 (.A(counter11_17_net_1), 
        .B(counter11_20_net_1), .C(counter11_19_net_1), .D(
        counter11_18_net_1), .Y(counter11_25_net_1));
    SLE \counter[12]  (.D(\counter_4[12]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[12]_net_1 ));
    SLE \counter[1]  (.D(un2_counter_1_cry_1_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[1]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \counter_4[21]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_21_S), .Y(\counter_4[21]_net_1 ));
    SLE \counter[3]  (.D(un2_counter_1_cry_3_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[3]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_7 (.A(VCC_net_1), .B(
        \counter[7]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_6_net_1), .S(un2_counter_1_cry_7_S), .Y(), 
        .FCO(un2_counter_1_cry_7_net_1));
    CFG2 #( .INIT(4'h4) )  \counter_4[17]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_17_S), .Y(\counter_4[17]_net_1 ));
    SLE \counter[23]  (.D(un2_counter_1_cry_23_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[23]_net_1 ));
    SLE \counter[19]  (.D(un2_counter_1_cry_19_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[19]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter11_20 (.A(\counter[31]_net_1 ), 
        .B(\counter[30]_net_1 ), .C(\counter[29]_net_1 ), .D(
        \counter[28]_net_1 ), .Y(counter11_20_net_1));
    CFG4 #( .INIT(16'h0001) )  counter12_17 (.A(\counter[15]_net_1 ), 
        .B(\counter[7]_net_1 ), .C(\counter[6]_net_1 ), .D(
        \counter[5]_net_1 ), .Y(counter12_17_net_1));
    CFG4 #( .INIT(16'h0001) )  counter11_19 (.A(\counter[27]_net_1 ), 
        .B(\counter[26]_net_1 ), .C(\counter[23]_net_1 ), .D(
        \counter[19]_net_1 ), .Y(counter11_19_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_23 (.A(VCC_net_1), 
        .B(\counter[23]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_22_net_1), .S(un2_counter_1_cry_23_S), .Y(), 
        .FCO(un2_counter_1_cry_23_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_2 (.A(VCC_net_1), .B(
        \counter[2]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_1_net_1), .S(un2_counter_1_cry_2_S), .Y(), 
        .FCO(un2_counter_1_cry_2_net_1));
    SLE \counter[20]  (.D(un2_counter_1_cry_20_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[20]_net_1 ));
    CFG2 #( .INIT(4'h4) )  \counter_4[12]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_12_S), .Y(\counter_4[12]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter12_16 (.A(\counter[4]_net_1 ), 
        .B(\counter[3]_net_1 ), .C(\counter[2]_net_1 ), .D(
        \counter[1]_net_1 ), .Y(counter12_16_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_17 (.A(VCC_net_1), 
        .B(\counter[17]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_16_net_1), .S(un2_counter_1_cry_17_S), .Y(), 
        .FCO(un2_counter_1_cry_17_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_6 (.A(VCC_net_1), .B(
        \counter[6]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_5_net_1), .S(un2_counter_1_cry_6_S), .Y(), 
        .FCO(un2_counter_1_cry_6_net_1));
    CFG4 #( .INIT(16'h8000) )  counter11_24 (.A(counter11_14_net_1), 
        .B(counter11_13_net_1), .C(counter11_16_net_1), .D(
        counter11_15_net_1), .Y(counter11_24_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_11 (.A(VCC_net_1), 
        .B(\counter[11]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_10_net_1), .S(un2_counter_1_cry_11_S), .Y(), 
        .FCO(un2_counter_1_cry_11_net_1));
    CFG2 #( .INIT(4'h1) )  \counter_4[0]  (.A(counter12_net_1), .B(
        \counter[0]_net_1 ), .Y(\counter_4[0]_net_1 ));
    SLE \counter[27]  (.D(un2_counter_1_cry_27_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[27]_net_1 ));
    SLE \counter[11]  (.D(\counter_4[11]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[11]_net_1 ));
    CFG4 #( .INIT(16'h0001) )  counter11_15 (.A(\counter[17]_net_1 ), 
        .B(\counter[14]_net_1 ), .C(\counter[12]_net_1 ), .D(
        \counter[9]_net_1 ), .Y(counter11_15_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_12 (.A(VCC_net_1), 
        .B(\counter[12]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_11_net_1), .S(un2_counter_1_cry_12_S), .Y(), 
        .FCO(un2_counter_1_cry_12_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_16 (.A(VCC_net_1), 
        .B(\counter[16]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_15_net_1), .S(un2_counter_1_cry_16_S), .Y(), 
        .FCO(un2_counter_1_cry_16_net_1));
    SLE \counter[30]  (.D(un2_counter_1_cry_30_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[30]_net_1 ));
    SLE \counter[18]  (.D(un2_counter_1_cry_18_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[18]_net_1 ));
    CFG4 #( .INIT(16'h8000) )  counter12_13 (.A(\counter[21]_net_1 ), 
        .B(\counter[17]_net_1 ), .C(\counter[14]_net_1 ), .D(
        \counter[12]_net_1 ), .Y(counter12_13_net_1));
    CFG2 #( .INIT(4'h4) )  \counter_4[14]  (.A(counter12_net_1), .B(
        un2_counter_1_cry_14_S), .Y(\counter_4[14]_net_1 ));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_25 (.A(VCC_net_1), 
        .B(\counter[25]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_24_net_1), .S(un2_counter_1_cry_25_S), .Y(), 
        .FCO(un2_counter_1_cry_25_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_30 (.A(VCC_net_1), 
        .B(\counter[30]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_29_net_1), .S(un2_counter_1_cry_30_S), .Y(), 
        .FCO(un2_counter_1_cry_30_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_24 (.A(VCC_net_1), 
        .B(\counter[24]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_23_net_1), .S(un2_counter_1_cry_24_S), .Y(), 
        .FCO(un2_counter_1_cry_24_net_1));
    CFG4 #( .INIT(16'h0001) )  counter12_18 (.A(\counter[27]_net_1 ), 
        .B(\counter[26]_net_1 ), .C(\counter[19]_net_1 ), .D(
        \counter[18]_net_1 ), .Y(counter12_18_net_1));
    CFG4 #( .INIT(16'h8000) )  counter11_14 (.A(\counter[24]_net_1 ), 
        .B(\counter[21]_net_1 ), .C(\counter[20]_net_1 ), .D(
        \counter[16]_net_1 ), .Y(counter11_14_net_1));
    CFG4 #( .INIT(16'h8000) )  counter12_24 (.A(counter12_18_net_1), 
        .B(counter12_17_net_1), .C(counter12_16_net_1), .D(
        counter11_20_net_1), .Y(counter12_24_net_1));
    ARI1 #( .INIT(20'h4AA00) )  un2_counter_1_cry_29 (.A(VCC_net_1), 
        .B(\counter[29]_net_1 ), .C(GND_net_1), .D(GND_net_1), .FCI(
        un2_counter_1_cry_28_net_1), .S(un2_counter_1_cry_29_S), .Y(), 
        .FCO(un2_counter_1_cry_29_net_1));
    SLE \counter[26]  (.D(un2_counter_1_cry_26_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[26]_net_1 ));
    SLE \counter[13]  (.D(un2_counter_1_cry_13_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[13]_net_1 ));
    SLE \counter[0]  (.D(\counter_4[0]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[0]_net_1 ));
    SLE \counter[10]  (.D(un2_counter_1_cry_10_S), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[10]_net_1 ));
    SLE \counter[9]  (.D(\counter_4[9]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[9]_net_1 ));
    SLE \counter[25]  (.D(\counter_4[25]_net_1 ), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(demo_0_MSS_READY), 
        .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(\counter[25]_net_1 ));
    
endmodule


module demo_FABOSC_0_OSC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC
    );
output FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;

    wire GND_net_1, VCC_net_1;
    
    RCOSC_25_50MHZ #( .FREQUENCY(50.0) )  I_RCOSC_25_50MHZ (.CLKOUT(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    
endmodule


module CoreResetP_Z1(
       demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N,
       demo_MSS_TMP_0_MSS_RESET_N_M2F,
       demo_0_POWER_ON_RESET_N,
       demo_0_FAB_CCC_GL0,
       demo_0_MSS_READY
    );
input  demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N;
input  demo_MSS_TMP_0_MSS_RESET_N_M2F;
input  demo_0_POWER_ON_RESET_N;
input  demo_0_FAB_CCC_GL0;
output demo_0_MSS_READY;

    wire MSS_HPMS_READY_int_net_1, mss_ready_select_net_1, VCC_net_1, 
        POWER_ON_RESET_N_clk_base_net_1, mss_ready_select4_net_1, 
        GND_net_1, mss_ready_state_net_1, RESET_N_M2F_clk_base_net_1, 
        POWER_ON_RESET_N_q1_net_1, RESET_N_M2F_q1_net_1, 
        FIC_2_APB_M_PRESET_N_clk_base_net_1, 
        FIC_2_APB_M_PRESET_N_q1_net_1, MSS_HPMS_READY_int_4_net_1;
    
    SLE RESET_N_M2F_clk_base (.D(RESET_N_M2F_q1_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        RESET_N_M2F_clk_base_net_1));
    SLE POWER_ON_RESET_N_clk_base (.D(POWER_ON_RESET_N_q1_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), .SLn(VCC_net_1), 
        .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_clk_base_net_1));
    SLE mss_ready_select (.D(VCC_net_1), .CLK(demo_0_FAB_CCC_GL0), .EN(
        mss_ready_select4_net_1), .ALn(POWER_ON_RESET_N_clk_base_net_1)
        , .ADn(VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(
        GND_net_1), .Q(mss_ready_select_net_1));
    CLKINT MSS_HPMS_READY_int_RNI3D75 (.A(MSS_HPMS_READY_int_net_1), 
        .Y(demo_0_MSS_READY));
    GND GND (.Y(GND_net_1));
    SLE mss_ready_state (.D(VCC_net_1), .CLK(demo_0_FAB_CCC_GL0), .EN(
        RESET_N_M2F_clk_base_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        mss_ready_state_net_1));
    VCC VCC (.Y(VCC_net_1));
    SLE RESET_N_M2F_q1 (.D(VCC_net_1), .CLK(demo_0_FAB_CCC_GL0), .EN(
        VCC_net_1), .ALn(demo_MSS_TMP_0_MSS_RESET_N_M2F), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(RESET_N_M2F_q1_net_1));
    SLE FIC_2_APB_M_PRESET_N_clk_base (.D(
        FIC_2_APB_M_PRESET_N_q1_net_1), .CLK(demo_0_FAB_CCC_GL0), .EN(
        VCC_net_1), .ALn(demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(
        VCC_net_1), .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), 
        .Q(FIC_2_APB_M_PRESET_N_clk_base_net_1));
    SLE POWER_ON_RESET_N_q1 (.D(VCC_net_1), .CLK(demo_0_FAB_CCC_GL0), 
        .EN(VCC_net_1), .ALn(demo_0_POWER_ON_RESET_N), .ADn(VCC_net_1), 
        .SLn(VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        POWER_ON_RESET_N_q1_net_1));
    CFG2 #( .INIT(4'h8) )  mss_ready_select4 (.A(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .B(mss_ready_state_net_1)
        , .Y(mss_ready_select4_net_1));
    CFG3 #( .INIT(8'hE0) )  MSS_HPMS_READY_int_4 (.A(
        RESET_N_M2F_clk_base_net_1), .B(mss_ready_select_net_1), .C(
        FIC_2_APB_M_PRESET_N_clk_base_net_1), .Y(
        MSS_HPMS_READY_int_4_net_1));
    SLE FIC_2_APB_M_PRESET_N_q1 (.D(VCC_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        FIC_2_APB_M_PRESET_N_q1_net_1));
    SLE MSS_HPMS_READY_int (.D(MSS_HPMS_READY_int_4_net_1), .CLK(
        demo_0_FAB_CCC_GL0), .EN(VCC_net_1), .ALn(
        POWER_ON_RESET_N_clk_base_net_1), .ADn(VCC_net_1), .SLn(
        VCC_net_1), .SD(GND_net_1), .LAT(GND_net_1), .Q(
        MSS_HPMS_READY_int_net_1));
    
endmodule


module demo_MSS(
       demo_0_FAB_CCC_GL0,
       LOCK,
       demo_MSS_TMP_0_MSS_RESET_N_M2F,
       demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N,
       MMUART_1_RXD,
       MMUART_1_TXD
    );
input  demo_0_FAB_CCC_GL0;
input  LOCK;
output demo_MSS_TMP_0_MSS_RESET_N_M2F;
output demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N;
input  MMUART_1_RXD;
output MMUART_1_TXD;

    wire MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT, 
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE, 
        MMUART_1_RXD_PAD_Y, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    MSS_075 #( .INIT(1438'h00000000000000000000000000000036100080000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000F00000000F000000000000000000000000000000007FFFFFFFB000001007C33F00000000E09500700003FFFFE400000000000010000000000F01C000001FE5FA4010842108421000001FE34001FF8000000400000000000451007FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF)
        , .ACT_UBITS(56'hFFFFFFFFFFFFFF), .MEMORYFILE("ENVM_init.mem")
        , .RTC_MAIN_XTL_FREQ(0.0), .RTC_MAIN_XTL_MODE(""), .DDR_CLK_FREQ(50.0)
         )  MSS_ADLIB_INST (.CAN_RXBUS_MGPIO3A_H2F_A(), 
        .CAN_RXBUS_MGPIO3A_H2F_B(), .CAN_TX_EBL_MGPIO4A_H2F_A(), 
        .CAN_TX_EBL_MGPIO4A_H2F_B(), .CAN_TXBUS_MGPIO2A_H2F_A(), 
        .CAN_TXBUS_MGPIO2A_H2F_B(), .CLK_CONFIG_APB(), .COMMS_INT(), 
        .CONFIG_PRESET_N(demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .EDAC_ERROR({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), 
        .F_FM0_RDATA({nc8, nc9, nc10, nc11, nc12, nc13, nc14, nc15, 
        nc16, nc17, nc18, nc19, nc20, nc21, nc22, nc23, nc24, nc25, 
        nc26, nc27, nc28, nc29, nc30, nc31, nc32, nc33, nc34, nc35, 
        nc36, nc37, nc38, nc39}), .F_FM0_READYOUT(), .F_FM0_RESP(), 
        .F_HM0_ADDR({nc40, nc41, nc42, nc43, nc44, nc45, nc46, nc47, 
        nc48, nc49, nc50, nc51, nc52, nc53, nc54, nc55, nc56, nc57, 
        nc58, nc59, nc60, nc61, nc62, nc63, nc64, nc65, nc66, nc67, 
        nc68, nc69, nc70, nc71}), .F_HM0_ENABLE(), .F_HM0_SEL(), 
        .F_HM0_SIZE({nc72, nc73}), .F_HM0_TRANS1(), .F_HM0_WDATA({nc74, 
        nc75, nc76, nc77, nc78, nc79, nc80, nc81, nc82, nc83, nc84, 
        nc85, nc86, nc87, nc88, nc89, nc90, nc91, nc92, nc93, nc94, 
        nc95, nc96, nc97, nc98, nc99, nc100, nc101, nc102, nc103, 
        nc104, nc105}), .F_HM0_WRITE(), .FAB_CHRGVBUS(), 
        .FAB_DISCHRGVBUS(), .FAB_DMPULLDOWN(), .FAB_DPPULLDOWN(), 
        .FAB_DRVVBUS(), .FAB_IDPULLUP(), .FAB_OPMODE({nc106, nc107}), 
        .FAB_SUSPENDM(), .FAB_TERMSEL(), .FAB_TXVALID(), .FAB_VCONTROL({
        nc108, nc109, nc110, nc111}), .FAB_VCONTROLLOADM(), 
        .FAB_XCVRSEL({nc112, nc113}), .FAB_XDATAOUT({nc114, nc115, 
        nc116, nc117, nc118, nc119, nc120, nc121}), .FACC_GLMUX_SEL(), 
        .FIC32_0_MASTER({nc122, nc123}), .FIC32_1_MASTER({nc124, nc125})
        , .FPGA_RESET_N(demo_MSS_TMP_0_MSS_RESET_N_M2F), .GTX_CLK(), 
        .H2F_INTERRUPT({nc126, nc127, nc128, nc129, nc130, nc131, 
        nc132, nc133, nc134, nc135, nc136, nc137, nc138, nc139, nc140, 
        nc141}), .H2F_NMI(), .H2FCALIB(), .I2C0_SCL_MGPIO31B_H2F_A(), 
        .I2C0_SCL_MGPIO31B_H2F_B(), .I2C0_SDA_MGPIO30B_H2F_A(), 
        .I2C0_SDA_MGPIO30B_H2F_B(), .I2C1_SCL_MGPIO1A_H2F_A(), 
        .I2C1_SCL_MGPIO1A_H2F_B(), .I2C1_SDA_MGPIO0A_H2F_A(), 
        .I2C1_SDA_MGPIO0A_H2F_B(), .MDCF(), .MDOENF(), .MDOF(), 
        .MMUART0_CTS_MGPIO19B_H2F_A(), .MMUART0_CTS_MGPIO19B_H2F_B(), 
        .MMUART0_DCD_MGPIO22B_H2F_A(), .MMUART0_DCD_MGPIO22B_H2F_B(), 
        .MMUART0_DSR_MGPIO20B_H2F_A(), .MMUART0_DSR_MGPIO20B_H2F_B(), 
        .MMUART0_DTR_MGPIO18B_H2F_A(), .MMUART0_DTR_MGPIO18B_H2F_B(), 
        .MMUART0_RI_MGPIO21B_H2F_A(), .MMUART0_RI_MGPIO21B_H2F_B(), 
        .MMUART0_RTS_MGPIO17B_H2F_A(), .MMUART0_RTS_MGPIO17B_H2F_B(), 
        .MMUART0_RXD_MGPIO28B_H2F_A(), .MMUART0_RXD_MGPIO28B_H2F_B(), 
        .MMUART0_SCK_MGPIO29B_H2F_A(), .MMUART0_SCK_MGPIO29B_H2F_B(), 
        .MMUART0_TXD_MGPIO27B_H2F_A(), .MMUART0_TXD_MGPIO27B_H2F_B(), 
        .MMUART1_DTR_MGPIO12B_H2F_A(), .MMUART1_RTS_MGPIO11B_H2F_A(), 
        .MMUART1_RTS_MGPIO11B_H2F_B(), .MMUART1_RXD_MGPIO26B_H2F_A(), 
        .MMUART1_RXD_MGPIO26B_H2F_B(), .MMUART1_SCK_MGPIO25B_H2F_A(), 
        .MMUART1_SCK_MGPIO25B_H2F_B(), .MMUART1_TXD_MGPIO24B_H2F_A(), 
        .MMUART1_TXD_MGPIO24B_H2F_B(), .MPLL_LOCK(), 
        .PER2_FABRIC_PADDR({nc142, nc143, nc144, nc145, nc146, nc147, 
        nc148, nc149, nc150, nc151, nc152, nc153, nc154, nc155}), 
        .PER2_FABRIC_PENABLE(), .PER2_FABRIC_PSEL(), 
        .PER2_FABRIC_PWDATA({nc156, nc157, nc158, nc159, nc160, nc161, 
        nc162, nc163, nc164, nc165, nc166, nc167, nc168, nc169, nc170, 
        nc171, nc172, nc173, nc174, nc175, nc176, nc177, nc178, nc179, 
        nc180, nc181, nc182, nc183, nc184, nc185, nc186, nc187}), 
        .PER2_FABRIC_PWRITE(), .RTC_MATCH(), .SLEEPDEEP(), 
        .SLEEPHOLDACK(), .SLEEPING(), .SMBALERT_NO0(), .SMBALERT_NO1(), 
        .SMBSUS_NO0(), .SMBSUS_NO1(), .SPI0_CLK_OUT(), 
        .SPI0_SDI_MGPIO5A_H2F_A(), .SPI0_SDI_MGPIO5A_H2F_B(), 
        .SPI0_SDO_MGPIO6A_H2F_A(), .SPI0_SDO_MGPIO6A_H2F_B(), 
        .SPI0_SS0_MGPIO7A_H2F_A(), .SPI0_SS0_MGPIO7A_H2F_B(), 
        .SPI0_SS1_MGPIO8A_H2F_A(), .SPI0_SS1_MGPIO8A_H2F_B(), 
        .SPI0_SS2_MGPIO9A_H2F_A(), .SPI0_SS2_MGPIO9A_H2F_B(), 
        .SPI0_SS3_MGPIO10A_H2F_A(), .SPI0_SS3_MGPIO10A_H2F_B(), 
        .SPI0_SS4_MGPIO19A_H2F_A(), .SPI0_SS5_MGPIO20A_H2F_A(), 
        .SPI0_SS6_MGPIO21A_H2F_A(), .SPI0_SS7_MGPIO22A_H2F_A(), 
        .SPI1_CLK_OUT(), .SPI1_SDI_MGPIO11A_H2F_A(), 
        .SPI1_SDI_MGPIO11A_H2F_B(), .SPI1_SDO_MGPIO12A_H2F_A(), 
        .SPI1_SDO_MGPIO12A_H2F_B(), .SPI1_SS0_MGPIO13A_H2F_A(), 
        .SPI1_SS0_MGPIO13A_H2F_B(), .SPI1_SS1_MGPIO14A_H2F_A(), 
        .SPI1_SS1_MGPIO14A_H2F_B(), .SPI1_SS2_MGPIO15A_H2F_A(), 
        .SPI1_SS2_MGPIO15A_H2F_B(), .SPI1_SS3_MGPIO16A_H2F_A(), 
        .SPI1_SS3_MGPIO16A_H2F_B(), .SPI1_SS4_MGPIO17A_H2F_A(), 
        .SPI1_SS5_MGPIO18A_H2F_A(), .SPI1_SS6_MGPIO23A_H2F_A(), 
        .SPI1_SS7_MGPIO24A_H2F_A(), .TCGF({nc188, nc189, nc190, nc191, 
        nc192, nc193, nc194, nc195, nc196, nc197}), .TRACECLK(), 
        .TRACEDATA({nc198, nc199, nc200, nc201}), .TX_CLK(), .TX_ENF(), 
        .TX_ERRF(), .TXCTL_EN_RIF(), .TXD_RIF({nc202, nc203, nc204, 
        nc205}), .TXDF({nc206, nc207, nc208, nc209, nc210, nc211, 
        nc212, nc213}), .TXEV(), .WDOGTIMEOUT(), .F_ARREADY_HREADYOUT1(
        ), .F_AWREADY_HREADYOUT0(), .F_BID({nc214, nc215, nc216, nc217})
        , .F_BRESP_HRESP0({nc218, nc219}), .F_BVALID(), 
        .F_RDATA_HRDATA01({nc220, nc221, nc222, nc223, nc224, nc225, 
        nc226, nc227, nc228, nc229, nc230, nc231, nc232, nc233, nc234, 
        nc235, nc236, nc237, nc238, nc239, nc240, nc241, nc242, nc243, 
        nc244, nc245, nc246, nc247, nc248, nc249, nc250, nc251, nc252, 
        nc253, nc254, nc255, nc256, nc257, nc258, nc259, nc260, nc261, 
        nc262, nc263, nc264, nc265, nc266, nc267, nc268, nc269, nc270, 
        nc271, nc272, nc273, nc274, nc275, nc276, nc277, nc278, nc279, 
        nc280, nc281, nc282, nc283}), .F_RID({nc284, nc285, nc286, 
        nc287}), .F_RLAST(), .F_RRESP_HRESP1({nc288, nc289}), 
        .F_RVALID(), .F_WREADY(), .MDDR_FABRIC_PRDATA({nc290, nc291, 
        nc292, nc293, nc294, nc295, nc296, nc297, nc298, nc299, nc300, 
        nc301, nc302, nc303, nc304, nc305}), .MDDR_FABRIC_PREADY(), 
        .MDDR_FABRIC_PSLVERR(), .CAN_RXBUS_F2H_SCP(VCC_net_1), 
        .CAN_TX_EBL_F2H_SCP(VCC_net_1), .CAN_TXBUS_F2H_SCP(VCC_net_1), 
        .COLF(VCC_net_1), .CRSF(VCC_net_1), .F2_DMAREADY({VCC_net_1, 
        VCC_net_1}), .F2H_INTERRUPT({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F2HCALIB(VCC_net_1), 
        .F_DMAREADY({VCC_net_1, VCC_net_1}), .F_FM0_ADDR({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_FM0_ENABLE(GND_net_1), .F_FM0_MASTLOCK(
        GND_net_1), .F_FM0_READY(VCC_net_1), .F_FM0_SEL(GND_net_1), 
        .F_FM0_SIZE({GND_net_1, GND_net_1}), .F_FM0_TRANS1(GND_net_1), 
        .F_FM0_WDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F_FM0_WRITE(GND_net_1), 
        .F_HM0_RDATA({GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1}), .F_HM0_READY(VCC_net_1), 
        .F_HM0_RESP(GND_net_1), .FAB_AVALID(VCC_net_1), 
        .FAB_HOSTDISCON(VCC_net_1), .FAB_IDDIG(VCC_net_1), 
        .FAB_LINESTATE({VCC_net_1, VCC_net_1}), .FAB_M3_RESET_N(
        VCC_net_1), .FAB_PLL_LOCK(LOCK), .FAB_RXACTIVE(VCC_net_1), 
        .FAB_RXERROR(VCC_net_1), .FAB_RXVALID(VCC_net_1), 
        .FAB_RXVALIDH(GND_net_1), .FAB_SESSEND(VCC_net_1), 
        .FAB_TXREADY(VCC_net_1), .FAB_VBUSVALID(VCC_net_1), 
        .FAB_VSTATUS({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), .FAB_XDATAIN({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .GTX_CLKPF(VCC_net_1), 
        .I2C0_BCLK(VCC_net_1), .I2C0_SCL_F2H_SCP(VCC_net_1), 
        .I2C0_SDA_F2H_SCP(VCC_net_1), .I2C1_BCLK(VCC_net_1), 
        .I2C1_SCL_F2H_SCP(VCC_net_1), .I2C1_SDA_F2H_SCP(VCC_net_1), 
        .MDIF(VCC_net_1), .MGPIO0A_F2H_GPIN(VCC_net_1), 
        .MGPIO10A_F2H_GPIN(VCC_net_1), .MGPIO11A_F2H_GPIN(VCC_net_1), 
        .MGPIO11B_F2H_GPIN(VCC_net_1), .MGPIO12A_F2H_GPIN(VCC_net_1), 
        .MGPIO13A_F2H_GPIN(VCC_net_1), .MGPIO14A_F2H_GPIN(VCC_net_1), 
        .MGPIO15A_F2H_GPIN(VCC_net_1), .MGPIO16A_F2H_GPIN(VCC_net_1), 
        .MGPIO17B_F2H_GPIN(VCC_net_1), .MGPIO18B_F2H_GPIN(VCC_net_1), 
        .MGPIO19B_F2H_GPIN(VCC_net_1), .MGPIO1A_F2H_GPIN(VCC_net_1), 
        .MGPIO20B_F2H_GPIN(VCC_net_1), .MGPIO21B_F2H_GPIN(VCC_net_1), 
        .MGPIO22B_F2H_GPIN(VCC_net_1), .MGPIO24B_F2H_GPIN(VCC_net_1), 
        .MGPIO25B_F2H_GPIN(VCC_net_1), .MGPIO26B_F2H_GPIN(VCC_net_1), 
        .MGPIO27B_F2H_GPIN(VCC_net_1), .MGPIO28B_F2H_GPIN(VCC_net_1), 
        .MGPIO29B_F2H_GPIN(VCC_net_1), .MGPIO2A_F2H_GPIN(VCC_net_1), 
        .MGPIO30B_F2H_GPIN(VCC_net_1), .MGPIO31B_F2H_GPIN(VCC_net_1), 
        .MGPIO3A_F2H_GPIN(VCC_net_1), .MGPIO4A_F2H_GPIN(VCC_net_1), 
        .MGPIO5A_F2H_GPIN(VCC_net_1), .MGPIO6A_F2H_GPIN(VCC_net_1), 
        .MGPIO7A_F2H_GPIN(VCC_net_1), .MGPIO8A_F2H_GPIN(VCC_net_1), 
        .MGPIO9A_F2H_GPIN(VCC_net_1), .MMUART0_CTS_F2H_SCP(VCC_net_1), 
        .MMUART0_DCD_F2H_SCP(VCC_net_1), .MMUART0_DSR_F2H_SCP(
        VCC_net_1), .MMUART0_DTR_F2H_SCP(VCC_net_1), 
        .MMUART0_RI_F2H_SCP(VCC_net_1), .MMUART0_RTS_F2H_SCP(VCC_net_1)
        , .MMUART0_RXD_F2H_SCP(VCC_net_1), .MMUART0_SCK_F2H_SCP(
        VCC_net_1), .MMUART0_TXD_F2H_SCP(VCC_net_1), 
        .MMUART1_CTS_F2H_SCP(VCC_net_1), .MMUART1_DCD_F2H_SCP(
        VCC_net_1), .MMUART1_DSR_F2H_SCP(VCC_net_1), 
        .MMUART1_RI_F2H_SCP(VCC_net_1), .MMUART1_RTS_F2H_SCP(VCC_net_1)
        , .MMUART1_RXD_F2H_SCP(VCC_net_1), .MMUART1_SCK_F2H_SCP(
        VCC_net_1), .MMUART1_TXD_F2H_SCP(VCC_net_1), 
        .PER2_FABRIC_PRDATA({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .PER2_FABRIC_PREADY(VCC_net_1), .PER2_FABRIC_PSLVERR(GND_net_1)
        , .RCGF({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .RX_CLKPF(VCC_net_1), .RX_DVF(VCC_net_1), .RX_ERRF(VCC_net_1), 
        .RX_EV(VCC_net_1), .RXDF({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .SLEEPHOLDREQ(GND_net_1), .SMBALERT_NI0(VCC_net_1), 
        .SMBALERT_NI1(VCC_net_1), .SMBSUS_NI0(VCC_net_1), .SMBSUS_NI1(
        VCC_net_1), .SPI0_CLK_IN(VCC_net_1), .SPI0_SDI_F2H_SCP(
        VCC_net_1), .SPI0_SDO_F2H_SCP(VCC_net_1), .SPI0_SS0_F2H_SCP(
        VCC_net_1), .SPI0_SS1_F2H_SCP(VCC_net_1), .SPI0_SS2_F2H_SCP(
        VCC_net_1), .SPI0_SS3_F2H_SCP(VCC_net_1), .SPI1_CLK_IN(
        VCC_net_1), .SPI1_SDI_F2H_SCP(VCC_net_1), .SPI1_SDO_F2H_SCP(
        VCC_net_1), .SPI1_SS0_F2H_SCP(VCC_net_1), .SPI1_SS1_F2H_SCP(
        VCC_net_1), .SPI1_SS2_F2H_SCP(VCC_net_1), .SPI1_SS3_F2H_SCP(
        VCC_net_1), .TX_CLKPF(VCC_net_1), .USER_MSS_GPIO_RESET_N(
        VCC_net_1), .USER_MSS_RESET_N(VCC_net_1), .XCLK_FAB(VCC_net_1), 
        .CLK_BASE(demo_0_FAB_CCC_GL0), .CLK_MDDR_APB(VCC_net_1), 
        .F_ARADDR_HADDR1({VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .F_ARBURST_HTRANS1({
        GND_net_1, GND_net_1}), .F_ARID_HSEL1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLEN_HBURST1({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_ARLOCK_HMASTLOCK1({GND_net_1, 
        GND_net_1}), .F_ARSIZE_HSIZE1({GND_net_1, GND_net_1}), 
        .F_ARVALID_HWRITE1(GND_net_1), .F_AWADDR_HADDR0({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_AWBURST_HTRANS0({GND_net_1, GND_net_1}), 
        .F_AWID_HSEL0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLEN_HBURST0({GND_net_1, GND_net_1, GND_net_1, GND_net_1}), 
        .F_AWLOCK_HMASTLOCK0({GND_net_1, GND_net_1}), .F_AWSIZE_HSIZE0({
        GND_net_1, GND_net_1}), .F_AWVALID_HWRITE0(GND_net_1), 
        .F_BREADY(GND_net_1), .F_RMW_AXI(GND_net_1), .F_RREADY(
        GND_net_1), .F_WDATA_HWDATA01({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .F_WID_HREADY01({GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .F_WLAST(GND_net_1), .F_WSTRB({GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1}), .F_WVALID(GND_net_1), 
        .FPGA_MDDR_ARESET_N(VCC_net_1), .MDDR_FABRIC_PADDR({VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1}), .MDDR_FABRIC_PENABLE(
        VCC_net_1), .MDDR_FABRIC_PSEL(VCC_net_1), .MDDR_FABRIC_PWDATA({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .MDDR_FABRIC_PWRITE(VCC_net_1), .PRESET_N(
        GND_net_1), .CAN_RXBUS_USBA_DATA1_MGPIO3A_IN(GND_net_1), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_IN(GND_net_1), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_IN(GND_net_1), .DM_IN({GND_net_1, 
        GND_net_1, GND_net_1}), .DRAM_DQ_IN({GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1, GND_net_1, GND_net_1, GND_net_1, GND_net_1, 
        GND_net_1}), .DRAM_DQS_IN({GND_net_1, GND_net_1, GND_net_1}), 
        .DRAM_FIFO_WE_IN({GND_net_1, GND_net_1}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_IN(GND_net_1), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_IN(GND_net_1), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_IN(GND_net_1), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_IN(GND_net_1), .MGPIO0B_IN(
        GND_net_1), .MGPIO10B_IN(GND_net_1), .MGPIO1B_IN(GND_net_1), 
        .MGPIO25A_IN(GND_net_1), .MGPIO26A_IN(GND_net_1), .MGPIO27A_IN(
        GND_net_1), .MGPIO28A_IN(GND_net_1), .MGPIO29A_IN(GND_net_1), 
        .MGPIO2B_IN(GND_net_1), .MGPIO30A_IN(GND_net_1), .MGPIO31A_IN(
        GND_net_1), .MGPIO3B_IN(GND_net_1), .MGPIO4B_IN(GND_net_1), 
        .MGPIO5B_IN(GND_net_1), .MGPIO6B_IN(GND_net_1), .MGPIO7B_IN(
        GND_net_1), .MGPIO8B_IN(GND_net_1), .MGPIO9B_IN(GND_net_1), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_IN(GND_net_1), 
        .MMUART0_DCD_MGPIO22B_IN(GND_net_1), .MMUART0_DSR_MGPIO20B_IN(
        GND_net_1), .MMUART0_DTR_USBC_DATA6_MGPIO18B_IN(GND_net_1), 
        .MMUART0_RI_MGPIO21B_IN(GND_net_1), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_IN(GND_net_1), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_IN(GND_net_1), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_IN(GND_net_1), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_IN(GND_net_1), 
        .MMUART1_CTS_MGPIO13B_IN(GND_net_1), .MMUART1_DCD_MGPIO16B_IN(
        GND_net_1), .MMUART1_DSR_MGPIO14B_IN(GND_net_1), 
        .MMUART1_DTR_MGPIO12B_IN(GND_net_1), .MMUART1_RI_MGPIO15B_IN(
        GND_net_1), .MMUART1_RTS_MGPIO11B_IN(GND_net_1), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_IN(MMUART_1_RXD_PAD_Y), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_IN(GND_net_1), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_IN(GND_net_1), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_IN(GND_net_1), 
        .RGMII_MDC_RMII_MDC_IN(GND_net_1), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_IN(GND_net_1), 
        .RGMII_RX_CLK_IN(GND_net_1), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_IN(GND_net_1), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_IN(GND_net_1), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_IN(GND_net_1), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_IN(GND_net_1), 
        .RGMII_RXD3_USBB_DATA4_IN(GND_net_1), .RGMII_TX_CLK_IN(
        GND_net_1), .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_IN(GND_net_1), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_IN(GND_net_1), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_IN(GND_net_1), 
        .RGMII_TXD2_USBB_DATA5_IN(GND_net_1), 
        .RGMII_TXD3_USBB_DATA6_IN(GND_net_1), .SPI0_SCK_USBA_XCLK_IN(
        GND_net_1), .SPI0_SDI_USBA_DIR_MGPIO5A_IN(GND_net_1), 
        .SPI0_SDO_USBA_STP_MGPIO6A_IN(GND_net_1), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_IN(GND_net_1), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_IN(GND_net_1), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_IN(GND_net_1), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_IN(GND_net_1), 
        .SPI0_SS4_MGPIO19A_IN(GND_net_1), .SPI0_SS5_MGPIO20A_IN(
        GND_net_1), .SPI0_SS6_MGPIO21A_IN(GND_net_1), 
        .SPI0_SS7_MGPIO22A_IN(GND_net_1), .SPI1_SCK_IN(GND_net_1), 
        .SPI1_SDI_MGPIO11A_IN(GND_net_1), .SPI1_SDO_MGPIO12A_IN(
        GND_net_1), .SPI1_SS0_MGPIO13A_IN(GND_net_1), 
        .SPI1_SS1_MGPIO14A_IN(GND_net_1), .SPI1_SS2_MGPIO15A_IN(
        GND_net_1), .SPI1_SS3_MGPIO16A_IN(GND_net_1), 
        .SPI1_SS4_MGPIO17A_IN(GND_net_1), .SPI1_SS5_MGPIO18A_IN(
        GND_net_1), .SPI1_SS6_MGPIO23A_IN(GND_net_1), 
        .SPI1_SS7_MGPIO24A_IN(GND_net_1), .USBC_XCLK_IN(GND_net_1), 
        .USBD_DATA0_IN(GND_net_1), .USBD_DATA1_IN(GND_net_1), 
        .USBD_DATA2_IN(GND_net_1), .USBD_DATA3_IN(GND_net_1), 
        .USBD_DATA4_IN(GND_net_1), .USBD_DATA5_IN(GND_net_1), 
        .USBD_DATA6_IN(GND_net_1), .USBD_DATA7_MGPIO23B_IN(GND_net_1), 
        .USBD_DIR_IN(GND_net_1), .USBD_NXT_IN(GND_net_1), .USBD_STP_IN(
        GND_net_1), .USBD_XCLK_IN(GND_net_1), 
        .CAN_RXBUS_USBA_DATA1_MGPIO3A_OUT(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OUT(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OUT(), .DRAM_ADDR({nc306, nc307, 
        nc308, nc309, nc310, nc311, nc312, nc313, nc314, nc315, nc316, 
        nc317, nc318, nc319, nc320, nc321}), .DRAM_BA({nc322, nc323, 
        nc324}), .DRAM_CASN(), .DRAM_CKE(), .DRAM_CLK(), .DRAM_CSN(), 
        .DRAM_DM_RDQS_OUT({nc325, nc326, nc327}), .DRAM_DQ_OUT({nc328, 
        nc329, nc330, nc331, nc332, nc333, nc334, nc335, nc336, nc337, 
        nc338, nc339, nc340, nc341, nc342, nc343, nc344, nc345}), 
        .DRAM_DQS_OUT({nc346, nc347, nc348}), .DRAM_FIFO_WE_OUT({nc349, 
        nc350}), .DRAM_ODT(), .DRAM_RASN(), .DRAM_RSTN(), .DRAM_WEN(), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OUT(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OUT(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OUT(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OUT(), .MGPIO0B_OUT(), 
        .MGPIO10B_OUT(), .MGPIO1B_OUT(), .MGPIO25A_OUT(), 
        .MGPIO26A_OUT(), .MGPIO27A_OUT(), .MGPIO28A_OUT(), 
        .MGPIO29A_OUT(), .MGPIO2B_OUT(), .MGPIO30A_OUT(), 
        .MGPIO31A_OUT(), .MGPIO3B_OUT(), .MGPIO4B_OUT(), .MGPIO5B_OUT()
        , .MGPIO6B_OUT(), .MGPIO7B_OUT(), .MGPIO8B_OUT(), .MGPIO9B_OUT(
        ), .MMUART0_CTS_USBC_DATA7_MGPIO19B_OUT(), 
        .MMUART0_DCD_MGPIO22B_OUT(), .MMUART0_DSR_MGPIO20B_OUT(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OUT(), 
        .MMUART0_RI_MGPIO21B_OUT(), 
        .MMUART0_RTS_USBC_DATA5_MGPIO17B_OUT(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OUT(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OUT(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OUT(), 
        .MMUART1_CTS_MGPIO13B_OUT(), .MMUART1_DCD_MGPIO16B_OUT(), 
        .MMUART1_DSR_MGPIO14B_OUT(), .MMUART1_DTR_MGPIO12B_OUT(), 
        .MMUART1_RI_MGPIO15B_OUT(), .MMUART1_RTS_MGPIO11B_OUT(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OUT(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OUT(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OUT(), 
        .RGMII_MDC_RMII_MDC_OUT(), 
        .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OUT(), .RGMII_RX_CLK_OUT(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OUT(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OUT(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OUT(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OUT(), 
        .RGMII_RXD3_USBB_DATA4_OUT(), .RGMII_TX_CLK_OUT(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OUT(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OUT(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OUT(), 
        .RGMII_TXD2_USBB_DATA5_OUT(), .RGMII_TXD3_USBB_DATA6_OUT(), 
        .SPI0_SCK_USBA_XCLK_OUT(), .SPI0_SDI_USBA_DIR_MGPIO5A_OUT(), 
        .SPI0_SDO_USBA_STP_MGPIO6A_OUT(), 
        .SPI0_SS0_USBA_NXT_MGPIO7A_OUT(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OUT(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OUT(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OUT(), .SPI0_SS4_MGPIO19A_OUT(), 
        .SPI0_SS5_MGPIO20A_OUT(), .SPI0_SS6_MGPIO21A_OUT(), 
        .SPI0_SS7_MGPIO22A_OUT(), .SPI1_SCK_OUT(), 
        .SPI1_SDI_MGPIO11A_OUT(), .SPI1_SDO_MGPIO12A_OUT(), 
        .SPI1_SS0_MGPIO13A_OUT(), .SPI1_SS1_MGPIO14A_OUT(), 
        .SPI1_SS2_MGPIO15A_OUT(), .SPI1_SS3_MGPIO16A_OUT(), 
        .SPI1_SS4_MGPIO17A_OUT(), .SPI1_SS5_MGPIO18A_OUT(), 
        .SPI1_SS6_MGPIO23A_OUT(), .SPI1_SS7_MGPIO24A_OUT(), 
        .USBC_XCLK_OUT(), .USBD_DATA0_OUT(), .USBD_DATA1_OUT(), 
        .USBD_DATA2_OUT(), .USBD_DATA3_OUT(), .USBD_DATA4_OUT(), 
        .USBD_DATA5_OUT(), .USBD_DATA6_OUT(), .USBD_DATA7_MGPIO23B_OUT(
        ), .USBD_DIR_OUT(), .USBD_NXT_OUT(), .USBD_STP_OUT(), 
        .USBD_XCLK_OUT(), .CAN_RXBUS_USBA_DATA1_MGPIO3A_OE(), 
        .CAN_TX_EBL_USBA_DATA2_MGPIO4A_OE(), 
        .CAN_TXBUS_USBA_DATA0_MGPIO2A_OE(), .DM_OE({nc351, nc352, 
        nc353}), .DRAM_DQ_OE({nc354, nc355, nc356, nc357, nc358, nc359, 
        nc360, nc361, nc362, nc363, nc364, nc365, nc366, nc367, nc368, 
        nc369, nc370, nc371}), .DRAM_DQS_OE({nc372, nc373, nc374}), 
        .I2C0_SCL_USBC_DATA1_MGPIO31B_OE(), 
        .I2C0_SDA_USBC_DATA0_MGPIO30B_OE(), 
        .I2C1_SCL_USBA_DATA4_MGPIO1A_OE(), 
        .I2C1_SDA_USBA_DATA3_MGPIO0A_OE(), .MGPIO0B_OE(), .MGPIO10B_OE(
        ), .MGPIO1B_OE(), .MGPIO25A_OE(), .MGPIO26A_OE(), .MGPIO27A_OE(
        ), .MGPIO28A_OE(), .MGPIO29A_OE(), .MGPIO2B_OE(), .MGPIO30A_OE(
        ), .MGPIO31A_OE(), .MGPIO3B_OE(), .MGPIO4B_OE(), .MGPIO5B_OE(), 
        .MGPIO6B_OE(), .MGPIO7B_OE(), .MGPIO8B_OE(), .MGPIO9B_OE(), 
        .MMUART0_CTS_USBC_DATA7_MGPIO19B_OE(), 
        .MMUART0_DCD_MGPIO22B_OE(), .MMUART0_DSR_MGPIO20B_OE(), 
        .MMUART0_DTR_USBC_DATA6_MGPIO18B_OE(), .MMUART0_RI_MGPIO21B_OE(
        ), .MMUART0_RTS_USBC_DATA5_MGPIO17B_OE(), 
        .MMUART0_RXD_USBC_STP_MGPIO28B_OE(), 
        .MMUART0_SCK_USBC_NXT_MGPIO29B_OE(), 
        .MMUART0_TXD_USBC_DIR_MGPIO27B_OE(), .MMUART1_CTS_MGPIO13B_OE()
        , .MMUART1_DCD_MGPIO16B_OE(), .MMUART1_DSR_MGPIO14B_OE(), 
        .MMUART1_DTR_MGPIO12B_OE(), .MMUART1_RI_MGPIO15B_OE(), 
        .MMUART1_RTS_MGPIO11B_OE(), 
        .MMUART1_RXD_USBC_DATA3_MGPIO26B_OE(), 
        .MMUART1_SCK_USBC_DATA4_MGPIO25B_OE(), 
        .MMUART1_TXD_USBC_DATA2_MGPIO24B_OE(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), 
        .RGMII_GTX_CLK_RMII_CLK_USBB_XCLK_OE(), .RGMII_MDC_RMII_MDC_OE(
        ), .RGMII_MDIO_RMII_MDIO_USBB_DATA7_OE(), .RGMII_RX_CLK_OE(), 
        .RGMII_RX_CTL_RMII_CRS_DV_USBB_DATA2_OE(), 
        .RGMII_RXD0_RMII_RXD0_USBB_DATA0_OE(), 
        .RGMII_RXD1_RMII_RXD1_USBB_DATA1_OE(), 
        .RGMII_RXD2_RMII_RX_ER_USBB_DATA3_OE(), 
        .RGMII_RXD3_USBB_DATA4_OE(), .RGMII_TX_CLK_OE(), 
        .RGMII_TX_CTL_RMII_TX_EN_USBB_NXT_OE(), 
        .RGMII_TXD0_RMII_TXD0_USBB_DIR_OE(), 
        .RGMII_TXD1_RMII_TXD1_USBB_STP_OE(), .RGMII_TXD2_USBB_DATA5_OE(
        ), .RGMII_TXD3_USBB_DATA6_OE(), .SPI0_SCK_USBA_XCLK_OE(), 
        .SPI0_SDI_USBA_DIR_MGPIO5A_OE(), .SPI0_SDO_USBA_STP_MGPIO6A_OE(
        ), .SPI0_SS0_USBA_NXT_MGPIO7A_OE(), 
        .SPI0_SS1_USBA_DATA5_MGPIO8A_OE(), 
        .SPI0_SS2_USBA_DATA6_MGPIO9A_OE(), 
        .SPI0_SS3_USBA_DATA7_MGPIO10A_OE(), .SPI0_SS4_MGPIO19A_OE(), 
        .SPI0_SS5_MGPIO20A_OE(), .SPI0_SS6_MGPIO21A_OE(), 
        .SPI0_SS7_MGPIO22A_OE(), .SPI1_SCK_OE(), .SPI1_SDI_MGPIO11A_OE(
        ), .SPI1_SDO_MGPIO12A_OE(), .SPI1_SS0_MGPIO13A_OE(), 
        .SPI1_SS1_MGPIO14A_OE(), .SPI1_SS2_MGPIO15A_OE(), 
        .SPI1_SS3_MGPIO16A_OE(), .SPI1_SS4_MGPIO17A_OE(), 
        .SPI1_SS5_MGPIO18A_OE(), .SPI1_SS6_MGPIO23A_OE(), 
        .SPI1_SS7_MGPIO24A_OE(), .USBC_XCLK_OE(), .USBD_DATA0_OE(), 
        .USBD_DATA1_OE(), .USBD_DATA2_OE(), .USBD_DATA3_OE(), 
        .USBD_DATA4_OE(), .USBD_DATA5_OE(), .USBD_DATA6_OE(), 
        .USBD_DATA7_MGPIO23B_OE(), .USBD_DIR_OE(), .USBD_NXT_OE(), 
        .USBD_STP_OE(), .USBD_XCLK_OE());
    GND GND (.Y(GND_net_1));
    TRIBUFF MMUART_1_TXD_PAD (.D(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OUT), .E(
        MSS_ADLIB_INST_MMUART1_TXD_USBC_DATA2_MGPIO24B_OE), .PAD(
        MMUART_1_TXD));
    INBUF MMUART_1_RXD_PAD (.PAD(MMUART_1_RXD), .Y(MMUART_1_RXD_PAD_Y));
    
endmodule


module demo_CCC_0_FCCC(
       FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC,
       LOCK,
       demo_0_FAB_CCC_GL0
    );
input  FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC;
output LOCK;
output demo_0_FAB_CCC_GL0;

    wire GL0_net, VCC_net_1, GND_net_1;
    
    VCC VCC (.Y(VCC_net_1));
    GND GND (.Y(GND_net_1));
    CLKINT GL0_INST (.A(GL0_net), .Y(demo_0_FAB_CCC_GL0));
    CCC #( .INIT(210'h0000007FB8000044D74000318C6318C1F18C61EC0404040400301)
        , .VCOFREQUENCY(800.0) )  CCC_INST (.Y0(), .Y1(), .Y2(), .Y3(), 
        .PRDATA({nc0, nc1, nc2, nc3, nc4, nc5, nc6, nc7}), .LOCK(LOCK), 
        .BUSY(), .CLK0(VCC_net_1), .CLK1(VCC_net_1), .CLK2(VCC_net_1), 
        .CLK3(VCC_net_1), .NGMUX0_SEL(GND_net_1), .NGMUX1_SEL(
        GND_net_1), .NGMUX2_SEL(GND_net_1), .NGMUX3_SEL(GND_net_1), 
        .NGMUX0_HOLD_N(VCC_net_1), .NGMUX1_HOLD_N(VCC_net_1), 
        .NGMUX2_HOLD_N(VCC_net_1), .NGMUX3_HOLD_N(VCC_net_1), 
        .NGMUX0_ARST_N(VCC_net_1), .NGMUX1_ARST_N(VCC_net_1), 
        .NGMUX2_ARST_N(VCC_net_1), .NGMUX3_ARST_N(VCC_net_1), 
        .PLL_BYPASS_N(VCC_net_1), .PLL_ARST_N(VCC_net_1), 
        .PLL_POWERDOWN_N(VCC_net_1), .GPD0_ARST_N(VCC_net_1), 
        .GPD1_ARST_N(VCC_net_1), .GPD2_ARST_N(VCC_net_1), .GPD3_ARST_N(
        VCC_net_1), .PRESET_N(GND_net_1), .PCLK(VCC_net_1), .PSEL(
        VCC_net_1), .PENABLE(VCC_net_1), .PWRITE(VCC_net_1), .PADDR({
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1}), .PWDATA({VCC_net_1, VCC_net_1, VCC_net_1, 
        VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1, VCC_net_1}), 
        .CLK0_PAD(GND_net_1), .CLK1_PAD(GND_net_1), .CLK2_PAD(
        GND_net_1), .CLK3_PAD(GND_net_1), .GL0(GL0_net), .GL1(), .GL2()
        , .GL3(), .RCOSC_25_50MHZ(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), 
        .RCOSC_1MHZ(GND_net_1), .XTLOSC(GND_net_1));
    
endmodule


module demo(
       MMUART_1_TXD,
       MMUART_1_RXD,
       demo_0_MSS_READY,
       demo_0_FAB_CCC_GL0,
       DEVRST_N,
       demo_0_POWER_ON_RESET_N
    );
output MMUART_1_TXD;
input  MMUART_1_RXD;
output demo_0_MSS_READY;
output demo_0_FAB_CCC_GL0;
input  DEVRST_N;
output demo_0_POWER_ON_RESET_N;

    wire SYSRESET_POR_net_1, 
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC, LOCK, 
        demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N, 
        demo_MSS_TMP_0_MSS_RESET_N_M2F, GND_net_1, VCC_net_1;
    
    demo_FABOSC_0_OSC FABOSC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC));
    CoreResetP_Z1 CORERESETP_0 (.demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N), 
        .demo_MSS_TMP_0_MSS_RESET_N_M2F(demo_MSS_TMP_0_MSS_RESET_N_M2F)
        , .demo_0_POWER_ON_RESET_N(demo_0_POWER_ON_RESET_N), 
        .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0), .demo_0_MSS_READY(
        demo_0_MSS_READY));
    VCC VCC (.Y(VCC_net_1));
    CLKINT SYSRESET_POR_RNIKPN2 (.A(SYSRESET_POR_net_1), .Y(
        demo_0_POWER_ON_RESET_N));
    demo_MSS demo_MSS_0 (.demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0), 
        .LOCK(LOCK), .demo_MSS_TMP_0_MSS_RESET_N_M2F(
        demo_MSS_TMP_0_MSS_RESET_N_M2F), 
        .demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N(
        demo_MSS_TMP_0_FIC_2_APB_M_PRESET_N), .MMUART_1_RXD(
        MMUART_1_RXD), .MMUART_1_TXD(MMUART_1_TXD));
    demo_CCC_0_FCCC CCC_0 (
        .FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC(
        FABOSC_0_RCOSC_25_50MHZ_CCC_OUT_RCOSC_25_50MHZ_CCC), .LOCK(
        LOCK), .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0));
    GND GND (.Y(GND_net_1));
    SYSRESET SYSRESET_POR (.POWER_ON_RESET_N(SYSRESET_POR_net_1), 
        .DEVRST_N(DEVRST_N));
    
endmodule


module demo_top(
       DEVRST_N,
       MMUART_1_RXD,
       LED1,
       LED2,
       LED3,
       LED4,
       MMUART_1_TXD
    );
input  DEVRST_N;
input  MMUART_1_RXD;
output LED1;
output LED2;
output LED3;
output LED4;
output MMUART_1_TXD;

    wire demo_0_FAB_CCC_GL0, demo_0_MSS_READY, demo_0_POWER_ON_RESET_N, 
        VCC_net_1, GND_net_1, LED1_c;
    
    OUTBUF LED4_obuf (.D(LED1_c), .PAD(LED4));
    OUTBUF LED1_obuf (.D(LED1_c), .PAD(LED1));
    Dev_Restart_after_ISP_blk Dev_Restart_after_ISP_blk_0 (
        .demo_0_POWER_ON_RESET_N(demo_0_POWER_ON_RESET_N), 
        .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0));
    VCC VCC (.Y(VCC_net_1));
    OUTBUF LED3_obuf (.D(LED1_c), .PAD(LED3));
    OUTBUF LED2_obuf (.D(LED1_c), .PAD(LED2));
    GND GND (.Y(GND_net_1));
    BLINK_LED BLINK_LED_0 (.LED1_c(LED1_c), .demo_0_FAB_CCC_GL0(
        demo_0_FAB_CCC_GL0), .demo_0_MSS_READY(demo_0_MSS_READY));
    demo demo_0 (.MMUART_1_TXD(MMUART_1_TXD), .MMUART_1_RXD(
        MMUART_1_RXD), .demo_0_MSS_READY(demo_0_MSS_READY), 
        .demo_0_FAB_CCC_GL0(demo_0_FAB_CCC_GL0), .DEVRST_N(DEVRST_N), 
        .demo_0_POWER_ON_RESET_N(demo_0_POWER_ON_RESET_N));
    
endmodule
