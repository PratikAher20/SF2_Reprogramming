`timescale 1 ns/100 ps
// Version: v11.5 11.5.0.26


module Dev_Restart_after_ISP_blk_TAMPER2_0_TAMPER2(
       RESET_N,
       JTAG_ACTIVE,
       LOCK_TAMPER_DETECT,
       MESH_SHORT_ERROR,
       DETECT_CATEGORY,
       DETECT_ATTEMPT,
       DETECT_FAIL,
       DIGEST_ERROR,
       SC_ROM_DIGEST_ERROR,
       TAMPER_CHANGE_STROBE
    );
input  RESET_N;
output JTAG_ACTIVE;
output LOCK_TAMPER_DETECT;
output MESH_SHORT_ERROR;
output [3:0] DETECT_CATEGORY;
output DETECT_ATTEMPT;
output DETECT_FAIL;
output DIGEST_ERROR;
output SC_ROM_DIGEST_ERROR;
output TAMPER_CHANGE_STROBE;

    wire VCC_NET;
    
    VCC VCC_INST (.Y(VCC_NET));
    TAMPER TAMPER_INST (.JTAG_ACTIVE(JTAG_ACTIVE), .LOCK_TAMPER_DETECT(
        LOCK_TAMPER_DETECT), .MESH_SHORT_ERROR(MESH_SHORT_ERROR), 
        .CLK_ERROR(), .DETECT_CATEGORY({DETECT_CATEGORY[3], 
        DETECT_CATEGORY[2], DETECT_CATEGORY[1], DETECT_CATEGORY[0]}), 
        .DETECT_ATTEMPT(DETECT_ATTEMPT), .DETECT_FAIL(DETECT_FAIL), 
        .DIGEST_ERROR(DIGEST_ERROR), .POWERUP_DIGEST_ERROR(), 
        .SC_ROM_DIGEST_ERROR(SC_ROM_DIGEST_ERROR), 
        .TAMPER_CHANGE_STROBE(TAMPER_CHANGE_STROBE), .LOCKDOWN_ALL_N(
        VCC_NET), .DISABLE_ALL_IOS_N(VCC_NET), .RESET_N(RESET_N), 
        .ZEROIZE_N(VCC_NET));
    
endmodule
